//
// Copyright (c) 2009-2017 Micron Technology, Inc. All Rights Reserved.
// This source code contains confidential information and trade secrets of
// Micron Technology, Inc.  Use, disclosure, or reproduction is prohibited
// without the prior express written permission of Micron Technology, Inc.
//
//

// *********************************************************
// UserWrapper
// This module instantiates the user module and all the stream and PicoBus
// connectors it needs.
//
// Macro defs:
//     PICOBUS_WIDTH       : enable pico bus
//     USER_MODULE_NAME    : enable user module, MUST have!
//     ENABLE_HMC          : enable hmc controller
//     ENABLE_2ND_HMC_LINK : enable 2nd hmc link (controller)
//     ENABLE_3RD_HMC_LINK : enable 3rd hmc link (controller)
//     ENABLE_4TH_HMC_LINK : enable 4th hmc link (controller)
//     USE_512_BIT_HMC_CONTROLLER : use the 1x512+1x128 port hmc controller, else use 5x128
//     ENABLE_QSPI_FLASH   : enable the quad SPI flash controller

//     STREAM*_IN_WIDTH    : enable * input stream
//     STREAM*_OUT_WIDTH   : enable * output stream
//
// *********************************************************

`include "PicoDefines.v"

module UserWrapper
    #(
`ifdef ENABLE_HMC
    parameter C_NUM_LINK                = 4 ,
`endif

`ifdef PICO_DDR3_OR_DDR4
`ifdef ALTERA_FPGA
    parameter AVL_DATA_WIDTH            = 512,
`ifdef PICO_DDR3
    parameter AVL_SIZE_WIDTH            = 9,
`elsif PICO_DDR4
    parameter AVL_SIZE_WIDTH            = 7,
`endif	// PICO_DDR
`ifdef PICO_MODEL_M506
    parameter AVL_ADDR_WIDTH            = 27,
`elsif PICO_MODEL_M520
    parameter AVL_ADDR_WIDTH            = 28,
`elsif PICO_MODEL_EX800
    parameter AVL_ADDR_WIDTH            = 26,
`endif	// PICO_MODEL
`endif	// ALTERA_FPGA
`ifdef PICO_MODEL_SB852
    parameter  ROW_WIDTH             =  17 ,
                                        // # of memory Row Address bits.
    parameter  CKE_WIDTH             =   2 ,
                                        // # of CKE outputs to memory.
    parameter  ODT_WIDTH             =   2 ,
                                        // # of ODT outputs to memory.
    parameter  DQ_WIDTH              =  72 ,
                                        // # of DQ (data)
    `ifdef SB852_16G
    parameter  DQS_WIDTH             =   9 ,
                                        // # of DQS/DQS# bits.
                                        // Number of DQS groups in I/O column #2.
    parameter  DBI_WIDTH             =   9 ,
    `else
    parameter  DQS_WIDTH             =  18 ,
                                        // 32G, 64G, 128G
    `ifdef SB852_64G
    parameter  CID_WIDTH             =   1 ,
    `elsif SB852_128G
    parameter  CID_WIDTH             =   2 ,
    `endif
    `endif
    parameter  CK_WIDTH              =   1 ,
                                        // # of CK/CK# outputs to memory.
    parameter nCS_PER_RANK              = 1,
                                        // # of unique CS outputs per Rank for
                                        // phy.
    parameter BANK_WIDTH                = 2,
`endif
            parameter C0_C_S_AXI_ID_WIDTH       = 12,   // width of the ID out of this UserWrapper
                                                        // = width of the ID from the masters + 4
            parameter C0_C_S_AXI_ADDR_WIDTH     = 32,   // AXI address width in MIG 0
            parameter C0_C_S_AXI_DATA_WIDTH     = 256,  // AXI data width in the MIG and interconnect
            parameter C0_C_S_AXI_MASTERS        = 3,    // number of master devices accessing MIG 0
`endif // PICO_DDR3_OR_DDR4
    parameter C_DATA_WIDTH		= 128,
    parameter OW_DVLD_W = (C_DATA_WIDTH==256)?'d2:'d1,
    parameter S_PB_RATIO = 62
    )

    (
`ifdef ENABLE_HMC
    input  wire                         hmc_tx_clk,
    input  wire                         hmc_rx_clk,
    input  wire                         hmc_rst,
    input  wire                         hmc_trained,

  `ifdef USE_512_BIT_HMC_CONTROLLER
    hmc_user_if                         hmc_port     [C_NUM_LINK-1:0] ,
    hmc_axi_if                          hmc_axi_port [C_NUM_LINK-1:0] ,

  `else //USE_512_BIT_HMC_CONTROLLER
    hmc_user_if                         hmc_port     [19:0] ,
  `endif //USE_512_BIT_HMC_CONTROLLER
    output wire                         PicoClk,
    output wire                         PicoRst,
    output wire [31:0]                  PicoAddr,
    output wire [`PICOBUS_WIDTH-1:0]    PicoDataIn,
    input  wire [`PICOBUS_WIDTH-1:0]    PicoDataOut,
    output wire                         PicoRd,
    output wire                         PicoWr,
`endif // ENABLE_HMC

`ifdef PICO_DDR3_OR_DDR4

        `ifdef PICO_MODEL_SB852
            input  wire                                c0_sys_clk_n    ,
            input  wire                                c0_sys_clk_p    ,
            input  wire                                c0_sys_rst_n    ,
            output wire                                c0_ddr4_act_n   ,
            output wire [ROW_WIDTH-1:0]                c0_ddr4_adr     ,
            output wire [BANK_WIDTH-1:0]               c0_ddr4_ba      ,
            output wire [BANK_WIDTH-1:0]               c0_ddr4_bg      ,
            output wire [CK_WIDTH-1:0]                 c0_ddr4_ck_c    ,
            output wire [CK_WIDTH-1:0]                 c0_ddr4_ck_t    ,
            output wire [CKE_WIDTH-1:0]                c0_ddr4_cke     ,
            output wire [BANK_WIDTH*nCS_PER_RANK-1:0]  c0_ddr4_cs_n    ,
            `ifdef SB852_16G
            inout  wire [DBI_WIDTH-1:0]                c0_ddr4_dm_n    ,
            `endif
            `ifdef SB852_64G
            output wire [CID_WIDTH-1:0]                c0_ddr4_c_id    ,
            `endif
            `ifdef SB852_128G
            output wire [CID_WIDTH-1:0]                c0_ddr4_c_id    ,
            `endif
            inout  wire [DQ_WIDTH-1:0]                 c0_ddr4_dq      ,
            inout  wire [DQS_WIDTH-1:0]                c0_ddr4_dqs_c   ,
            inout  wire [DQS_WIDTH-1:0]                c0_ddr4_dqs_t   ,
            output wire [ODT_WIDTH-1:0]                c0_ddr4_odt     ,
            output wire                                c0_ddr4_par     ,
            output wire                                c0_ddr4_reset_n ,

            input  wire                                c1_sys_clk_n    ,
            input  wire                                c1_sys_clk_p    ,
            input  wire                                c1_sys_rst_n    ,
            output wire                                c1_ddr4_act_n   ,
            output wire [ROW_WIDTH-1:0]                c1_ddr4_adr     ,
            output wire [BANK_WIDTH-1:0]               c1_ddr4_ba      ,
            output wire [BANK_WIDTH-1:0]               c1_ddr4_bg      ,
            output wire [CK_WIDTH-1:0]                 c1_ddr4_ck_c    ,
            output wire [CK_WIDTH-1:0]                 c1_ddr4_ck_t    ,
            output wire [CKE_WIDTH-1:0]                c1_ddr4_cke     ,
            output wire [BANK_WIDTH*nCS_PER_RANK-1:0]  c1_ddr4_cs_n    ,
            `ifdef SB852_16G
            inout  wire [DBI_WIDTH-1:0]                c1_ddr4_dm_n    ,
            `endif
            `ifdef SB852_64G
            output wire [CID_WIDTH-1:0]                c1_ddr4_c_id    ,
            `endif
            `ifdef SB852_128G
            output wire [CID_WIDTH-1:0]                c1_ddr4_c_id    ,
            `endif
            inout  wire [DQ_WIDTH-1:0]                 c1_ddr4_dq      ,
            inout  wire [DQS_WIDTH-1:0]                c1_ddr4_dqs_c   ,
            inout  wire [DQS_WIDTH-1:0]                c1_ddr4_dqs_t   ,
            output wire [ODT_WIDTH-1:0]                c1_ddr4_odt     ,
            output wire                                c1_ddr4_par     ,
            output wire                                c1_ddr4_reset_n ,

            input  wire                                c2_sys_clk_n    ,
            input  wire                                c2_sys_clk_p    ,
            input  wire                                c2_sys_rst_n    ,
            output wire                                c2_ddr4_act_n   ,
            output wire [ROW_WIDTH-1:0]                c2_ddr4_adr     ,
            output wire [BANK_WIDTH-1:0]               c2_ddr4_ba      ,
            output wire [BANK_WIDTH-1:0]               c2_ddr4_bg      ,
            output wire [CK_WIDTH-1:0]                 c2_ddr4_ck_c    ,
            output wire [CK_WIDTH-1:0]                 c2_ddr4_ck_t    ,
            output wire [CKE_WIDTH-1:0]                c2_ddr4_cke     ,
            output wire [BANK_WIDTH*nCS_PER_RANK-1:0]  c2_ddr4_cs_n    ,
            `ifdef SB852_16G
            inout  wire [DBI_WIDTH-1:0]                c2_ddr4_dm_n    ,
            `endif
            `ifdef SB852_64G
            output wire [CID_WIDTH-1:0]                c2_ddr4_c_id    ,
            `endif
            `ifdef SB852_128G
            output wire [CID_WIDTH-1:0]                c2_ddr4_c_id    ,
            `endif
            inout  wire [DQ_WIDTH-1:0]                 c2_ddr4_dq      ,
            inout  wire [DQS_WIDTH-1:0]                c2_ddr4_dqs_c   ,
            inout  wire [DQS_WIDTH-1:0]                c2_ddr4_dqs_t   ,
            output wire [ODT_WIDTH-1:0]                c2_ddr4_odt     ,
            output wire                                c2_ddr4_par     ,
            output wire                                c2_ddr4_reset_n ,

            input  wire                                c3_sys_clk_n    ,
            input  wire                                c3_sys_clk_p    ,
            input  wire                                c3_sys_rst_n    ,
            output wire                                c3_ddr4_act_n   ,
            output wire [ROW_WIDTH-1:0]                c3_ddr4_adr     ,
            output wire [BANK_WIDTH-1:0]               c3_ddr4_ba      ,
            output wire [BANK_WIDTH-1:0]               c3_ddr4_bg      ,
            output wire [CK_WIDTH-1:0]                 c3_ddr4_ck_c    ,
            output wire [CK_WIDTH-1:0]                 c3_ddr4_ck_t    ,
            output wire [CKE_WIDTH-1:0]                c3_ddr4_cke     ,
            output wire [BANK_WIDTH*nCS_PER_RANK-1:0]  c3_ddr4_cs_n    ,
            `ifdef SB852_16G
            inout  wire [DBI_WIDTH-1:0]                c3_ddr4_dm_n    ,
            `endif
            `ifdef SB852_64G
            output wire [CID_WIDTH-1:0]                c3_ddr4_c_id    ,
            `endif
            `ifdef SB852_128G
            output wire [CID_WIDTH-1:0]                c3_ddr4_c_id    ,
            `endif
            inout  wire [DQ_WIDTH-1:0]                 c3_ddr4_dq      ,
            inout  wire [DQS_WIDTH-1:0]                c3_ddr4_dqs_c   ,
            inout  wire [DQS_WIDTH-1:0]                c3_ddr4_dqs_t   ,
            output wire [ODT_WIDTH-1:0]                c3_ddr4_odt     ,
            output wire                                c3_ddr4_par     ,
            output wire                                c3_ddr4_reset_n ,
    `else
	    //------------------------------------------------------
	    // DDR3 Reset
	    //------------------------------------------------------
        output [0:0]                         ddr3_sys_rst,        // Resets the DDR3
    `endif

	//------------------------------------------------------
	// DDR3 0  - AXI ports
	//------------------------------------------------------
      input                                c0_tb_clk,           // AXI input clock

      // Input control signals
      `ifndef PICO_MODEL_SB852
          input                                c0_phy_init_done,    // Initialization completed
      `endif
      input                                c0_tb_rst,           // Active high reset signal
`ifdef ALTERA_FPGA
    input  wire                                 avl_ready,
    output wire   [AVL_ADDR_WIDTH-1:0]          avl_addr,
    input  wire                                 avl_rdata_valid,
    input  wire   [AVL_DATA_WIDTH-1:0]          avl_rdata,
    output wire   [AVL_DATA_WIDTH-1:0]          avl_wdata,
    output wire   [AVL_DATA_WIDTH/8-1:0]        avl_be,
    output wire                                 avl_read_req,
    output wire                                 avl_write_req,
    output wire   [AVL_SIZE_WIDTH-1:0]          avl_size,
`else
      // AXI write address channel signals
      input                                c0_s_axi_awready,    // Indicates slave is ready to accept a
      output [C0_C_S_AXI_ID_WIDTH-1:0]     c0_s_axi_awid,       // Write ID
      output [C0_C_S_AXI_ADDR_WIDTH-1:0]   c0_s_axi_awaddr,     // Write address
      output [7:0]                         c0_s_axi_awlen,      // Write Burst Length
      output [2:0]                         c0_s_axi_awsize,     // Write Burst size
      output [1:0]                         c0_s_axi_awburst,    // Write Burst type
      output                               c0_s_axi_awlock,     // Write lock type
      output [3:0]                         c0_s_axi_awcache,    // Write Cache type
      output [2:0]                         c0_s_axi_awprot,     // Write Protection type
      output [3:0]                         c0_s_axi_awqos,      // Write Quality of Service Signaling
      output                               c0_s_axi_awvalid,    // Write address valid

      // AXI write data channel signals
      input                                c0_s_axi_wready,     // Write data ready
      output [C0_C_S_AXI_DATA_WIDTH-1:0]   c0_s_axi_wdata,      // Write data
      output [C0_C_S_AXI_DATA_WIDTH/8-1:0] c0_s_axi_wstrb,      // Write strobes
      output                               c0_s_axi_wlast,      // Last write transaction
      output                               c0_s_axi_wvalid,     // Write valid

      // AXI write response channel signals
      input  [C0_C_S_AXI_ID_WIDTH-1:0]     c0_s_axi_bid,        // Response ID
      input  [1:0]                         c0_s_axi_bresp,      // Write response
      input                                c0_s_axi_bvalid,     // Write reponse valid
      output                               c0_s_axi_bready,     // Response ready

      // AXI read address channel signals
      input                                c0_s_axi_arready,    // Read address ready
      output [C0_C_S_AXI_ID_WIDTH-1:0]     c0_s_axi_arid,       // Read ID
      output [C0_C_S_AXI_ADDR_WIDTH-1:0]   c0_s_axi_araddr,     // Read address
      output [7:0]                         c0_s_axi_arlen,      // Read Burst Length
      output [2:0]                         c0_s_axi_arsize,     // Read Burst size
      output [1:0]                         c0_s_axi_arburst,    // Read Burst type
      output                               c0_s_axi_arlock,     // Read lock type
      output [3:0]                         c0_s_axi_arcache,    // Read Cache type
      output [2:0]                         c0_s_axi_arprot,     // Read Protection type
      output                               c0_s_axi_arvalid,    // Read address valid
      output [3:0]                         c0_s_axi_arqos,      // Read Quality of Service Signaling

      // AXI read data channel signals
      input  [C0_C_S_AXI_ID_WIDTH-1:0]     c0_s_axi_rid,        // Response ID
      input  [1:0]                         c0_s_axi_rresp,      // Read response
      input                                c0_s_axi_rvalid,     // Read reponse valid
      input  [C0_C_S_AXI_DATA_WIDTH-1:0]   c0_s_axi_rdata,      // Read data
      input                                c0_s_axi_rlast,      // Read last
      output                               c0_s_axi_rready,     // Read Response ready

`endif // ALTERA_FPGA
`endif // PICO_DDR3_OR_DDR4

    input               extra_clk,
    input               clk,
    input               rst,

`ifdef USER_DIRECT_PCI
    // user-direct writes
    output [C_DATA_WIDTH-1:0]      user_pci_wr_q_data,
    output              user_pci_wr_q_valid,
    input               user_pci_wr_q_en,

    output [C_DATA_WIDTH-1:0]      user_pci_wr_data_q_data,
    output              user_pci_wr_data_q_valid,
    input               user_pci_wr_data_q_en,

    input               direct_rx_valid,
`endif // USER_DIRECT_PCI

    input  [OW_DVLD_W-1:0] s_out_en,
    input  [8:0]        s_out_id,
    output [C_DATA_WIDTH-1:0] s_out_data,
    output [OW_DVLD_W-1:0] s_out_ow_dvld,

    input               s_in_valid,
    input [8:0]         s_in_id,
    input [C_DATA_WIDTH-1:0] s_in_data,
    input [OW_DVLD_W-1:0] s_in_ow_dvld,

    input       [8:0]   s_poll_id,
    output      [31:0]  s_poll_seq,
    output      [127:0] s_poll_next_desc,
    output              s_poll_next_desc_valid,

    input       [8:0]   s_next_desc_rd_id,
    input               s_next_desc_rd_en

// Add the I2C pins to connect to the CPLD on the SB852
`ifdef PICO_MODEL_SB852
  `ifdef ENABLE_QSPI_FLASH
    ,
    inout               scl,
    inout               sda
  `endif
`endif



    );

    // function to compute ceil( log( x ) )
    // Note: log is computed in base 2
    function integer clogb2;
        input [31:0] value;
        begin
            value = value - 1;
            for (clogb2 = 0; value > 0; clogb2 = clogb2 + 1) begin
                value = value >> 1;
            end
        end
    endfunction

    `ifdef USER_MODULE_NAME                 // Only enable these streams if there is a usermodule

    /////////////////////////////////
    // UserModule PicoBus
    /////////////////////////////////
`ifdef PICOBUS_WIDTH
        wire [C_DATA_WIDTH-1:0] s_out_data_userpb;
	wire [OW_DVLD_W-1:0] s_out_ow_dvld_userpb;
	wire [127:0]    s_poll_next_desc_userpb;
        wire [31:0]     s_poll_seq_userpb;
        wire            s_poll_next_desc_valid_userpb;

        wire [`PICOBUS_WIDTH-1:0]   UserModulePicoDataIn, UserModulePicoDataOut;
        wire [31:0]                 UserModulePicoAddr;
        wire                        UserModulePicoClk, UserModulePicoRst, UserModulePicoRd, UserModulePicoWr;
`endif // PICOBUS_WIDTH

    wire [31:0]     stream_in_desc_poll_seq[127:0];
    wire            stream_in_desc_poll_next_desc_valid[127:0];
    wire [127:0]    stream_in_desc_poll_next_desc[127:0];

    wire            stream_in_rdy[127:0];
    wire            stream_in_valid[127:0];
    wire [C_DATA_WIDTH-1:0] stream_in_data[127:0];
    wire [OW_DVLD_W-1:0] stream_in_ow_dvld[127:0];

    wire [31:0]     stream_out_desc_poll_seq[127:0];
    wire            stream_out_desc_poll_next_desc_valid[127:0];
    wire [127:0]    stream_out_desc_poll_next_desc[127:0];
    wire [C_DATA_WIDTH-1:0] stream_out_data_card[127:0];        // This has to be ored together
    wire [OW_DVLD_W-1:0] stream_out_ow_dvld_card[127:0];        // This has to be ored together

    wire            stream_out_rdy[127:0];
    wire            stream_out_valid[127:0];
    wire [C_DATA_WIDTH-1:0] stream_out_data[127:0];
    wire [OW_DVLD_W-1:0] stream_out_ow_dvld[127:0];

    //////////////////////////////
    // STREAM TO Flash Controller
    //////////////////////////////

`ifdef ENABLE_QSPI_FLASH
    // QSPI flash controller for the SB852 and optionally other Xilinx based modules
    // Connected via 128-bit output stream ID 115 and input stream ID 115

    StreamToFlashCtl #( .WIDTH      (64),        // PicoBus width
                        .S_PB_RATIO (2)          // 250MHz stream clock, 125 MHz flash_ctl clk, 62.5MHz SPI clock
                      ) StreamToFlashCtl (
                        .s_clk             (clk),
                        .s_rst             (rst),

                        .si_ready          (stream_in_rdy[`FLASH_CTL_STREAM_ID]),
                        .si_valid          (stream_in_valid[`FLASH_CTL_STREAM_ID]),
                        .si_data           (stream_in_data[`FLASH_CTL_STREAM_ID][127:0]),

                        .so_ready          (stream_out_rdy[`FLASH_CTL_STREAM_ID]),
                        .so_valid          (stream_out_valid[`FLASH_CTL_STREAM_ID]),
                        .so_data           (stream_out_data[`FLASH_CTL_STREAM_ID][127:0]),

                        .scl               (scl),
                        .sda               (sda)

                      );
`endif // ENABLE_QSPI_FLASH

    ///////////////////
    // STREAM TO HMC
    ///////////////////

`ifdef ENABLE_HMC
    // Note: we assume that if the HMC is being used, then PICOBUS_WIDTH has
    // defined to be 32.
    assign PicoClk          = UserModulePicoClk;
    assign PicoRst          = UserModulePicoRst;
    assign PicoRd           = UserModulePicoRd;
    assign PicoWr           = UserModulePicoWr;
    assign PicoAddr         = UserModulePicoAddr;
    assign PicoDataIn       = UserModulePicoDataIn;

    // stream to HMC port[0]
    PicoStreamToHMC #(
        .C_AXI_ID_WIDTH     (6),
        .C_AXI_ADDR_WIDTH   (34),
        .C_AXI_DATA_WIDTH   (128)
    )
    stream_to_hmc_0
    (
        // streaming interface
        .clk                (clk),
        .rst                (rst),

        .si_ready           (stream_in_rdy[`HMC_STREAM_ID]),
        .si_valid           (stream_in_valid[`HMC_STREAM_ID]),
        .si_data            (stream_in_data[`HMC_STREAM_ID][127:0]),
        .so_ready           (stream_out_rdy[`HMC_STREAM_ID]),
        .so_valid           (stream_out_valid[`HMC_STREAM_ID]),
        .so_data            (stream_out_data[`HMC_STREAM_ID][127:0]),

        // HMC port signals
        .hmc_tx_clk                         (hmc_tx_clk),
        .hmc_rx_clk                         (hmc_rx_clk),
        .hmc_rst                            (hmc_rst),
        .hmc_trained                        (hmc_trained),

        .hmc_clk                            ( hmc_port[0].clk ),
        .hmc_addr                           ( hmc_port[0].addr ),
        .hmc_size                           ( hmc_port[0].size ),
        .hmc_tag                            ( hmc_port[0].tag ),
        .hmc_cmd_valid                      ( hmc_port[0].cmd_valid ),
        .hmc_cmd_ready                      ( hmc_port[0].cmd_ready ),
        .hmc_cmd                            ( hmc_port[0].cmd ),
        .hmc_wr_data                        ( hmc_port[0].wr_data ),
        .hmc_wr_data_valid                  ( hmc_port[0].wr_data_valid ),
        .hmc_wr_data_ready                  ( hmc_port[0].wr_data_ready ),

        .hmc_rd_data                        ( hmc_port[0].rd_data ),
        .hmc_rd_data_tag                    ( hmc_port[0].rd_data_tag ),
        .hmc_rd_data_valid                  ( hmc_port[0].rd_data_valid ),
        .hmc_errstat                        ( hmc_port[0].errstat ),
        .hmc_dinv                           ( hmc_port[0].dinv )
    );
`endif // ENABLE_HMC


`ifdef PICO_DDR3_OR_DDR4

    ////////////////
    // DDR3 MIG 0 //
    ////////////////
    // Slave Interface Wires
    wire    [C0_C_S_AXI_MASTERS:0]          c0_axi_clk;

    // Slave Interface Write Address Ports
    wire    [C0_C_S_AXI_ID_WIDTH-5:0]       c0_axi_awid    [0:C0_C_S_AXI_MASTERS];
    wire    [C0_C_S_AXI_ADDR_WIDTH-1:0]     c0_axi_awaddr  [0:C0_C_S_AXI_MASTERS];
    wire    [7:0]                           c0_axi_awlen   [0:C0_C_S_AXI_MASTERS];
    wire    [2:0]                           c0_axi_awsize  [0:C0_C_S_AXI_MASTERS];
    wire    [1:0]                           c0_axi_awburst [0:C0_C_S_AXI_MASTERS];
    wire    [0:0]                           c0_axi_awlock  [0:C0_C_S_AXI_MASTERS];
    wire    [3:0]                           c0_axi_awcache [0:C0_C_S_AXI_MASTERS];
    wire    [2:0]                           c0_axi_awprot  [0:C0_C_S_AXI_MASTERS];
    wire    [3:0]                           c0_axi_awqos   [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_awvalid [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_awready [0:C0_C_S_AXI_MASTERS];
    // Slave Interface Write Data Ports
    wire    [C0_C_S_AXI_DATA_WIDTH-1:0]     c0_axi_wdata   [0:C0_C_S_AXI_MASTERS];
    wire    [C0_C_S_AXI_DATA_WIDTH/8-1:0]   c0_axi_wstrb   [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_wlast   [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_wvalid  [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_wready  [0:C0_C_S_AXI_MASTERS];
    // Slave Interface Write Response Ports
    wire    [C0_C_S_AXI_ID_WIDTH-5:0]       c0_axi_bid     [0:C0_C_S_AXI_MASTERS];
    wire    [1:0]                           c0_axi_bresp   [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_bvalid  [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_bready  [0:C0_C_S_AXI_MASTERS];
    // Slave Interface Read Address Ports
    wire    [C0_C_S_AXI_ID_WIDTH-5:0]       c0_axi_arid    [0:C0_C_S_AXI_MASTERS];
    wire    [C0_C_S_AXI_ADDR_WIDTH-1:0]     c0_axi_araddr  [0:C0_C_S_AXI_MASTERS];
    wire    [7:0]                           c0_axi_arlen   [0:C0_C_S_AXI_MASTERS];
    wire    [2:0]                           c0_axi_arsize  [0:C0_C_S_AXI_MASTERS];
    wire    [1:0]                           c0_axi_arburst [0:C0_C_S_AXI_MASTERS];
    wire    [0:0]                           c0_axi_arlock  [0:C0_C_S_AXI_MASTERS];
    wire    [3:0]                           c0_axi_arcache [0:C0_C_S_AXI_MASTERS];
    wire    [2:0]                           c0_axi_arprot  [0:C0_C_S_AXI_MASTERS];
    wire    [3:0]                           c0_axi_arqos   [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_arvalid [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_arready [0:C0_C_S_AXI_MASTERS];
    // Slave Interface Read Data Ports
    wire    [C0_C_S_AXI_ID_WIDTH-5:0]       c0_axi_rid     [0:C0_C_S_AXI_MASTERS];
    wire    [C0_C_S_AXI_DATA_WIDTH-1:0]     c0_axi_rdata   [0:C0_C_S_AXI_MASTERS];
    wire    [1:0]                           c0_axi_rresp   [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_rlast   [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_rvalid  [0:C0_C_S_AXI_MASTERS];
    wire                                    c0_axi_rready  [0:C0_C_S_AXI_MASTERS];

`ifdef PICO_MODEL_SB852
    wire   [0:0]                            ddr3_sys_rst;
    wire                                    c0_phy_init_done;
    wire                                    c0_clk;
    wire                                    c0_rst;
    wire                                    c1_clk;
    wire                                    c1_rst;
    wire                                    c2_clk;
    wire                                    c2_rst;
    wire                                    c3_clk;
    wire                                    c3_rst;

    mem_subsystem_wrapper #(

    ) PicoMemSubsytem (
    .S00_ACLK          ( clk                ),
    .S00_ARESETN       (~rst                ),
    .S00_AXI_araddr    ( c0_axi_araddr  [0] ),
    .S00_AXI_arburst   ( c0_axi_arburst [0] ),
    .S00_AXI_arcache   ( c0_axi_arcache [0] ),
    .S00_AXI_arid      ( c0_axi_arid    [0] ),
    .S00_AXI_arlen     ( c0_axi_arlen   [0] ),
    .S00_AXI_arlock    ( c0_axi_arlock  [0] ),
    .S00_AXI_arprot    ( c0_axi_arprot  [0] ),
    .S00_AXI_arqos     ( c0_axi_arqos   [0] ),
    .S00_AXI_arready   ( c0_axi_arready [0] ),
    .S00_AXI_arregion  ( 4'd0               ),
    .S00_AXI_arsize    ( c0_axi_arsize  [0] ),
    .S00_AXI_arvalid   ( c0_axi_arvalid [0] ),
    .S00_AXI_awaddr    ( c0_axi_awaddr  [0] ),
    .S00_AXI_awburst   ( c0_axi_awburst [0] ),
    .S00_AXI_awcache   ( c0_axi_awcache [0] ),
    .S00_AXI_awid      ( c0_axi_awid    [0] ),
    .S00_AXI_awlen     ( c0_axi_awlen   [0] ),
    .S00_AXI_awlock    ( c0_axi_awlock  [0] ),
    .S00_AXI_awprot    ( c0_axi_awprot  [0] ),
    .S00_AXI_awqos     ( c0_axi_awqos   [0] ),
    .S00_AXI_awready   ( c0_axi_awready [0] ),
    .S00_AXI_awregion  ( 4'd0               ),
    .S00_AXI_awsize    ( c0_axi_awsize  [0] ),
    .S00_AXI_awvalid   ( c0_axi_awvalid [0] ),
    .S00_AXI_bid       ( c0_axi_bid     [0] ),
    .S00_AXI_bready    ( c0_axi_bready  [0] ),
    .S00_AXI_bresp     ( c0_axi_bresp   [0] ),
    .S00_AXI_bvalid    ( c0_axi_bvalid  [0] ),
    .S00_AXI_rdata     ( c0_axi_rdata   [0] ),
    .S00_AXI_rid       ( c0_axi_rid     [0] ),
    .S00_AXI_rlast     ( c0_axi_rlast   [0] ),
    .S00_AXI_rready    ( c0_axi_rready  [0] ),
    .S00_AXI_rresp     ( c0_axi_rresp   [0] ),
    .S00_AXI_rvalid    ( c0_axi_rvalid  [0] ),
    .S00_AXI_wdata     ( c0_axi_wdata   [0] ),
    .S00_AXI_wlast     ( c0_axi_wlast   [0] ),
    .S00_AXI_wready    ( c0_axi_wready  [0] ),
    .S00_AXI_wstrb     ( c0_axi_wstrb   [0] ),
    .S00_AXI_wvalid    ( c0_axi_wvalid  [0] ),

    .S01_ACLK          ( c0_axi_clk     [1] ),
    .S01_ARESETN       (~c0_rst             ),
    .S01_AXI_araddr    ( c0_axi_araddr  [1] ),
    .S01_AXI_arburst   ( c0_axi_arburst [1] ),
    .S01_AXI_arcache   ( c0_axi_arcache [1] ),
    .S01_AXI_arid      ( c0_axi_arid    [1] ),
    .S01_AXI_arlen     ( c0_axi_arlen   [1] ),
    .S01_AXI_arlock    ( c0_axi_arlock  [1] ),
    .S01_AXI_arprot    ( c0_axi_arprot  [1] ),
    .S01_AXI_arqos     ( c0_axi_arqos   [1] ),
    .S01_AXI_arready   ( c0_axi_arready [1] ),
    .S01_AXI_arregion  ( 4'd0               ),
    .S01_AXI_arsize    ( c0_axi_arsize  [1] ),
    .S01_AXI_arvalid   ( c0_axi_arvalid [1] ),
    .S01_AXI_awaddr    ( c0_axi_awaddr  [1] ),
    .S01_AXI_awburst   ( c0_axi_awburst [1] ),
    .S01_AXI_awcache   ( c0_axi_awcache [1] ),
    .S01_AXI_awid      ( c0_axi_awid    [1] ),
    .S01_AXI_awlen     ( c0_axi_awlen   [1] ),
    .S01_AXI_awlock    ( c0_axi_awlock  [1] ),
    .S01_AXI_awprot    ( c0_axi_awprot  [1] ),
    .S01_AXI_awqos     ( c0_axi_awqos   [1] ),
    .S01_AXI_awready   ( c0_axi_awready [1] ),
    .S01_AXI_awregion  ( 4'd0               ),
    .S01_AXI_awsize    ( c0_axi_awsize  [1] ),
    .S01_AXI_awvalid   ( c0_axi_awvalid [1] ),
    .S01_AXI_bid       ( c0_axi_bid     [1] ),
    .S01_AXI_bready    ( c0_axi_bready  [1] ),
    .S01_AXI_bresp     ( c0_axi_bresp   [1] ),
    .S01_AXI_bvalid    ( c0_axi_bvalid  [1] ),
    .S01_AXI_rdata     ( c0_axi_rdata   [1] ),
    .S01_AXI_rid       ( c0_axi_rid     [1] ),
    .S01_AXI_rlast     ( c0_axi_rlast   [1] ),
    .S01_AXI_rready    ( c0_axi_rready  [1] ),
    .S01_AXI_rresp     ( c0_axi_rresp   [1] ),
    .S01_AXI_rvalid    ( c0_axi_rvalid  [1] ),
    .S01_AXI_wdata     ( c0_axi_wdata   [1] ),
    .S01_AXI_wlast     ( c0_axi_wlast   [1] ),
    .S01_AXI_wready    ( c0_axi_wready  [1] ),
    .S01_AXI_wstrb     ( c0_axi_wstrb   [1] ),
    .S01_AXI_wvalid    ( c0_axi_wvalid  [1] ),

    //.S02_ACLK          ( clk                ),
    //.S02_ARESETN       (~rst                ),
    //.S02_AXI_araddr    ( c0_axi_araddr  [2] ),
    //.S02_AXI_arburst   ( c0_axi_arburst [2] ),
    //.S02_AXI_arcache   ( c0_axi_arcache [2] ),
    //.S02_AXI_arid      ( c0_axi_arid    [2] ),
    //.S02_AXI_arlen     ( c0_axi_arlen   [2] ),
    //.S02_AXI_arlock    ( c0_axi_arlock  [2] ),
    //.S02_AXI_arprot    ( c0_axi_arprot  [2] ),
    //.S02_AXI_arqos     ( c0_axi_arqos   [2] ),
    //.S02_AXI_arready   ( c0_axi_arready [2] ),
    //.S02_AXI_arregion  ( 4'd0               ),
    //.S02_AXI_arsize    ( c0_axi_arsize  [2] ),
    //.S02_AXI_arvalid   ( c0_axi_arvalid [2] ),
    //.S02_AXI_awaddr    ( c0_axi_awaddr  [2] ),
    //.S02_AXI_awburst   ( c0_axi_awburst [2] ),
    //.S02_AXI_awcache   ( c0_axi_awcache [2] ),
    //.S02_AXI_awid      ( c0_axi_awid    [2] ),
    //.S02_AXI_awlen     ( c0_axi_awlen   [2] ),
    //.S02_AXI_awlock    ( c0_axi_awlock  [2] ),
    //.S02_AXI_awprot    ( c0_axi_awprot  [2] ),
    //.S02_AXI_awqos     ( c0_axi_awqos   [2] ),
    //.S02_AXI_awready   ( c0_axi_awready [2] ),
    //.S02_AXI_awregion  ( 4'd0               ),
    //.S02_AXI_awsize    ( c0_axi_awsize  [2] ),
    //.S02_AXI_awvalid   ( c0_axi_awvalid [2] ),
    //.S02_AXI_bid       ( c0_axi_bid     [2] ),
    //.S02_AXI_bready    ( c0_axi_bready  [2] ),
    //.S02_AXI_bresp     ( c0_axi_bresp   [2] ),
    //.S02_AXI_bvalid    ( c0_axi_bvalid  [2] ),
    //.S02_AXI_rdata     ( c0_axi_rdata   [2] ),
    //.S02_AXI_rid       ( c0_axi_rid     [2] ),
    //.S02_AXI_rlast     ( c0_axi_rlast   [2] ),
    //.S02_AXI_rready    ( c0_axi_rready  [2] ),
    //.S02_AXI_rresp     ( c0_axi_rresp   [2] ),
    //.S02_AXI_rvalid    ( c0_axi_rvalid  [2] ),
    //.S02_AXI_wdata     ( c0_axi_wdata   [2] ),
    //.S02_AXI_wlast     ( c0_axi_wlast   [2] ),
    //.S02_AXI_wready    ( c0_axi_wready  [2] ),
    //.S02_AXI_wstrb     ( c0_axi_wstrb   [2] ),
    //.S02_AXI_wvalid    ( c0_axi_wvalid  [2] ),

    //.S03_ACLK          ( clk                ),
    //.S03_ARESETN       (~rst                ),
    //.S03_AXI_araddr    ( c0_axi_araddr  [3] ),
    //.S03_AXI_arburst   ( c0_axi_arburst [3] ),
    //.S03_AXI_arcache   ( c0_axi_arcache [3] ),
    //.S03_AXI_arid      ( c0_axi_arid    [3] ),
    //.S03_AXI_arlen     ( c0_axi_arlen   [3] ),
    //.S03_AXI_arlock    ( c0_axi_arlock  [3] ),
    //.S03_AXI_arprot    ( c0_axi_arprot  [3] ),
    //.S03_AXI_arqos     ( c0_axi_arqos   [3] ),
    //.S03_AXI_arready   ( c0_axi_arready [3] ),
    //.S03_AXI_arregion  ( 4'd0               ),
    //.S03_AXI_arsize    ( c0_axi_arsize  [3] ),
    //.S03_AXI_arvalid   ( c0_axi_arvalid [3] ),
    //.S03_AXI_awaddr    ( c0_axi_awaddr  [3] ),
    //.S03_AXI_awburst   ( c0_axi_awburst [3] ),
    //.S03_AXI_awcache   ( c0_axi_awcache [3] ),
    //.S03_AXI_awid      ( c0_axi_awid    [3] ),
    //.S03_AXI_awlen     ( c0_axi_awlen   [3] ),
    //.S03_AXI_awlock    ( c0_axi_awlock  [3] ),
    //.S03_AXI_awprot    ( c0_axi_awprot  [3] ),
    //.S03_AXI_awqos     ( c0_axi_awqos   [3] ),
    //.S03_AXI_awready   ( c0_axi_awready [3] ),
    //.S03_AXI_awregion  ( 4'd0               ),
    //.S03_AXI_awsize    ( c0_axi_awsize  [3] ),
    //.S03_AXI_awvalid   ( c0_axi_awvalid [3] ),
    //.S03_AXI_bid       ( c0_axi_bid     [3] ),
    //.S03_AXI_bready    ( c0_axi_bready  [3] ),
    //.S03_AXI_bresp     ( c0_axi_bresp   [3] ),
    //.S03_AXI_bvalid    ( c0_axi_bvalid  [3] ),
    //.S03_AXI_rdata     ( c0_axi_rdata   [3] ),
    //.S03_AXI_rid       ( c0_axi_rid     [3] ),
    //.S03_AXI_rlast     ( c0_axi_rlast   [3] ),
    //.S03_AXI_rready    ( c0_axi_rready  [3] ),
    //.S03_AXI_rresp     ( c0_axi_rresp   [3] ),
    //.S03_AXI_rvalid    ( c0_axi_rvalid  [3] ),
    //.S03_AXI_wdata     ( c0_axi_wdata   [3] ),
    //.S03_AXI_wlast     ( c0_axi_wlast   [3] ),
    //.S03_AXI_wready    ( c0_axi_wready  [3] ),
    //.S03_AXI_wstrb     ( c0_axi_wstrb   [3] ),
    //.S03_AXI_wvalid    ( c0_axi_wvalid  [3] ),

    //.S04_ACLK          ( clk                ),
    //.S04_ARESETN       (~rst                ),
    //.S04_AXI_araddr    ( c0_axi_araddr  [4] ),
    //.S04_AXI_arburst   ( c0_axi_arburst [4] ),
    //.S04_AXI_arcache   ( c0_axi_arcache [4] ),
    //.S04_AXI_arid      ( c0_axi_arid    [4] ),
    //.S04_AXI_arlen     ( c0_axi_arlen   [4] ),
    //.S04_AXI_arlock    ( c0_axi_arlock  [4] ),
    //.S04_AXI_arprot    ( c0_axi_arprot  [4] ),
    //.S04_AXI_arqos     ( c0_axi_arqos   [4] ),
    //.S04_AXI_arready   ( c0_axi_arready [4] ),
    //.S04_AXI_arregion  ( 4'd0               ),
    //.S04_AXI_arsize    ( c0_axi_arsize  [4] ),
    //.S04_AXI_arvalid   ( c0_axi_arvalid [4] ),
    //.S04_AXI_awaddr    ( c0_axi_awaddr  [4] ),
    //.S04_AXI_awburst   ( c0_axi_awburst [4] ),
    //.S04_AXI_awcache   ( c0_axi_awcache [4] ),
    //.S04_AXI_awid      ( c0_axi_awid    [4] ),
    //.S04_AXI_awlen     ( c0_axi_awlen   [4] ),
    //.S04_AXI_awlock    ( c0_axi_awlock  [4] ),
    //.S04_AXI_awprot    ( c0_axi_awprot  [4] ),
    //.S04_AXI_awqos     ( c0_axi_awqos   [4] ),
    //.S04_AXI_awready   ( c0_axi_awready [4] ),
    //.S04_AXI_awregion  ( 4'd0               ),
    //.S04_AXI_awsize    ( c0_axi_awsize  [4] ),
    //.S04_AXI_awvalid   ( c0_axi_awvalid [4] ),
    //.S04_AXI_bid       ( c0_axi_bid     [4] ),
    //.S04_AXI_bready    ( c0_axi_bready  [4] ),
    //.S04_AXI_bresp     ( c0_axi_bresp   [4] ),
    //.S04_AXI_bvalid    ( c0_axi_bvalid  [4] ),
    //.S04_AXI_rdata     ( c0_axi_rdata   [4] ),
    //.S04_AXI_rid       ( c0_axi_rid     [4] ),
    //.S04_AXI_rlast     ( c0_axi_rlast   [4] ),
    //.S04_AXI_rready    ( c0_axi_rready  [4] ),
    //.S04_AXI_rresp     ( c0_axi_rresp   [4] ),
    //.S04_AXI_rvalid    ( c0_axi_rvalid  [4] ),
    //.S04_AXI_wdata     ( c0_axi_wdata   [4] ),
    //.S04_AXI_wlast     ( c0_axi_wlast   [4] ),
    //.S04_AXI_wready    ( c0_axi_wready  [4] ),
    //.S04_AXI_wstrb     ( c0_axi_wstrb   [4] ),
    //.S04_AXI_wvalid    ( c0_axi_wvalid  [4] ),

    .c0_clk            ( c0_clk             ),
    .c0_rst            ( c0_rst             ),

    .c0_sys_clk_n      ( c0_sys_clk_n       ),
    .c0_sys_clk_p      ( c0_sys_clk_p       ),
    .c0_sys_rst_n      ( c0_sys_rst_n & ~ddr3_sys_rst ),
    .c0_ddr4_act_n     ( c0_ddr4_act_n      ),
    .c0_ddr4_adr       ( c0_ddr4_adr        ),
    .c0_ddr4_ba        ( c0_ddr4_ba         ),
    .c0_ddr4_bg        ( c0_ddr4_bg         ),
    .c0_ddr4_ck_c      ( c0_ddr4_ck_c       ),
    .c0_ddr4_ck_t      ( c0_ddr4_ck_t       ),
    .c0_ddr4_cke       ( c0_ddr4_cke        ),
    .c0_ddr4_cs_n      ( c0_ddr4_cs_n       ),
    .c0_ddr4_dq        ( c0_ddr4_dq         ),
    .c0_ddr4_dqs_c     ( c0_ddr4_dqs_c      ),
    .c0_ddr4_dqs_t     ( c0_ddr4_dqs_t      ),
    .c0_ddr4_odt       ( c0_ddr4_odt        ),
    .c0_ddr4_par       ( c0_ddr4_par        ),
    .c0_ddr4_reset_n   ( c0_ddr4_reset_n    ),
    `ifdef SB852_16G
    .c0_ddr4_dm_n      ( c0_ddr4_dm_n       ),
    `endif
    `ifdef SB852_64G
    .c0_ddr4_c_id      ( c0_ddr4_c_id       ),
    `endif
    `ifdef SB852_128G
    .c0_ddr4_c_id      ( c0_ddr4_c_id       ),
    `endif
    
    .c1_clk            ( c1_clk             ),
    .c1_rst            ( c1_rst             ),

    .c1_sys_clk_n      ( c1_sys_clk_n       ),
    .c1_sys_clk_p      ( c1_sys_clk_p       ),
    .c1_sys_rst_n      ( c1_sys_rst_n & ~ddr3_sys_rst ),
    .c1_ddr4_act_n     ( c1_ddr4_act_n      ),
    .c1_ddr4_adr       ( c1_ddr4_adr        ),
    .c1_ddr4_ba        ( c1_ddr4_ba         ),
    .c1_ddr4_bg        ( c1_ddr4_bg         ),
    .c1_ddr4_ck_c      ( c1_ddr4_ck_c       ),
    .c1_ddr4_ck_t      ( c1_ddr4_ck_t       ),
    .c1_ddr4_cke       ( c1_ddr4_cke        ),
    .c1_ddr4_cs_n      ( c1_ddr4_cs_n       ),
    .c1_ddr4_dq        ( c1_ddr4_dq         ),
    .c1_ddr4_dqs_c     ( c1_ddr4_dqs_c      ),
    .c1_ddr4_dqs_t     ( c1_ddr4_dqs_t      ),
    .c1_ddr4_odt       ( c1_ddr4_odt        ),
    .c1_ddr4_par       ( c1_ddr4_par        ),
    .c1_ddr4_reset_n   ( c1_ddr4_reset_n    ),
    `ifdef SB852_16G
    .c1_ddr4_dm_n      ( c1_ddr4_dm_n       ),
    `endif
    `ifdef SB852_64G
    .c1_ddr4_c_id      ( c1_ddr4_c_id       ),
    `endif
    `ifdef SB852_128G
    .c1_ddr4_c_id      ( c1_ddr4_c_id       ),
    `endif
        
    .c2_clk            ( c2_clk             ),
    .c2_rst            ( c2_rst             ),

    .c2_sys_clk_n      ( c2_sys_clk_n       ),
    .c2_sys_clk_p      ( c2_sys_clk_p       ),
    .c2_sys_rst_n      ( c2_sys_rst_n & ~ddr3_sys_rst ),
    .c2_ddr4_act_n     ( c2_ddr4_act_n      ),
    .c2_ddr4_adr       ( c2_ddr4_adr        ),
    .c2_ddr4_ba        ( c2_ddr4_ba         ),
    .c2_ddr4_bg        ( c2_ddr4_bg         ),
    .c2_ddr4_ck_c      ( c2_ddr4_ck_c       ),
    .c2_ddr4_ck_t      ( c2_ddr4_ck_t       ),
    .c2_ddr4_cke       ( c2_ddr4_cke        ),
    .c2_ddr4_cs_n      ( c2_ddr4_cs_n       ),
    .c2_ddr4_dq        ( c2_ddr4_dq         ),
    .c2_ddr4_dqs_c     ( c2_ddr4_dqs_c      ),
    .c2_ddr4_dqs_t     ( c2_ddr4_dqs_t      ),
    .c2_ddr4_odt       ( c2_ddr4_odt        ),
    .c2_ddr4_par       ( c2_ddr4_par        ),
    .c2_ddr4_reset_n   ( c2_ddr4_reset_n    ),
    `ifdef SB852_16G
    .c2_ddr4_dm_n      ( c2_ddr4_dm_n       ),
    `endif
    `ifdef SB852_64G
    .c2_ddr4_c_id      ( c2_ddr4_c_id       ),
    `endif
    `ifdef SB852_128G
    .c2_ddr4_c_id      ( c2_ddr4_c_id       ),
    `endif
        
    .c3_clk            ( c3_clk             ),
    .c3_rst            ( c3_rst             ),

    .c3_sys_clk_n      ( c3_sys_clk_n       ),
    .c3_sys_clk_p      ( c3_sys_clk_p       ),
    .c3_sys_rst_n      ( c3_sys_rst_n & ~ddr3_sys_rst ),
    .c3_ddr4_act_n     ( c3_ddr4_act_n      ),
    .c3_ddr4_adr       ( c3_ddr4_adr        ),
    .c3_ddr4_ba        ( c3_ddr4_ba         ),
    .c3_ddr4_bg        ( c3_ddr4_bg         ),
    .c3_ddr4_ck_c      ( c3_ddr4_ck_c       ),
    .c3_ddr4_ck_t      ( c3_ddr4_ck_t       ),
    .c3_ddr4_cke       ( c3_ddr4_cke        ),
    .c3_ddr4_cs_n      ( c3_ddr4_cs_n       ),
    .c3_ddr4_dq        ( c3_ddr4_dq         ),
    .c3_ddr4_dqs_c     ( c3_ddr4_dqs_c      ),
    .c3_ddr4_dqs_t     ( c3_ddr4_dqs_t      ),
    .c3_ddr4_odt       ( c3_ddr4_odt        ),
    .c3_ddr4_par       ( c3_ddr4_par        ),
    .c3_ddr4_reset_n   ( c3_ddr4_reset_n    ),
    `ifdef SB852_16G
    .c3_ddr4_dm_n      ( c3_ddr4_dm_n       ),
    `endif
    `ifdef SB852_64G
    .c3_ddr4_c_id      ( c3_ddr4_c_id       ),
    `endif
    `ifdef SB852_128G
    .c3_ddr4_c_id      ( c3_ddr4_c_id       ),
    `endif
    .ddr_calib_complete( c0_phy_init_done   )
    );

`else

    PicoAXIInterconnect #(
`ifdef PICO_DDR4
    `ifdef ALTERA_FPGA
        // for altera different MEM size
        .AVL_ADDR_WIDTH         (AVL_ADDR_WIDTH),
        .AVL_DATA_WIDTH         (AVL_DATA_WIDTH),
        .AVL_SIZE_WIDTH         (AVL_SIZE_WIDTH),
    `endif
`endif // PICO_DDR4
        .PICO_AXI_MASTERS       (C0_C_S_AXI_MASTERS+1),
        .C_AXI_ID_WIDTH         (C0_C_S_AXI_ID_WIDTH),
        .C_AXI_ADDR_WIDTH       (C0_C_S_AXI_ADDR_WIDTH),
        .C_AXI_DATA_WIDTH       (C0_C_S_AXI_DATA_WIDTH)
    ) new_axi_ic (
        .ddr3_ui_clk        (c0_tb_clk),
        .ddr3_ui_rst        (c0_tb_rst),

        .clk                (clk),
        .rst                (rst),

        .s0_axi_clk         (c0_axi_clk[0]),
        .s0_axi_awid        (c0_axi_awid[0]),
        .s0_axi_awaddr      (c0_axi_awaddr[0]),
        .s0_axi_awlen       (c0_axi_awlen[0]),
        .s0_axi_awsize      (c0_axi_awsize[0]),
        .s0_axi_awburst     (c0_axi_awburst[0]),
        .s0_axi_awlock      (c0_axi_awlock[0]),
        .s0_axi_awcache     (c0_axi_awcache[0]),
        .s0_axi_awprot      (c0_axi_awprot[0]),
        .s0_axi_awqos       (c0_axi_awqos[0]),
        .s0_axi_awvalid     (c0_axi_awvalid[0]),
        .s0_axi_awready     (c0_axi_awready[0]),
        .s0_axi_wdata       (c0_axi_wdata[0]),
        .s0_axi_wstrb       (c0_axi_wstrb[0]),
        .s0_axi_wlast       (c0_axi_wlast[0]),
        .s0_axi_wvalid      (c0_axi_wvalid[0]),
        .s0_axi_wready      (c0_axi_wready[0]),
        .s0_axi_bid         (c0_axi_bid[0]),
        .s0_axi_bresp       (c0_axi_bresp[0]),
        .s0_axi_bvalid      (c0_axi_bvalid[0]),
        .s0_axi_bready      (c0_axi_bready[0]),
        .s0_axi_arid        (c0_axi_arid[0]),
        .s0_axi_araddr      (c0_axi_araddr[0]),
        .s0_axi_arlen       (c0_axi_arlen[0]),
        .s0_axi_arsize      (c0_axi_arsize[0]),
        .s0_axi_arburst     (c0_axi_arburst[0]),
        .s0_axi_arlock      (c0_axi_arlock[0]),
        .s0_axi_arcache     (c0_axi_arcache[0]),
        .s0_axi_arprot      (c0_axi_arprot[0]),
        .s0_axi_arqos       (c0_axi_arqos[0]),
        .s0_axi_arvalid     (c0_axi_arvalid[0]),
        .s0_axi_arready     (c0_axi_arready[0]),
        .s0_axi_rid         (c0_axi_rid[0]),
        .s0_axi_rdata       (c0_axi_rdata[0]),
        .s0_axi_rresp       (c0_axi_rresp[0]),
        .s0_axi_rlast       (c0_axi_rlast[0]),
        .s0_axi_rvalid      (c0_axi_rvalid[0]),
        .s0_axi_rready      (c0_axi_rready[0]),

   `ifdef PICO_AXI_PORT_1
        // master port 1
        .s1_axi_clk      (c0_axi_clk[1]),
        .s1_axi_awid     (c0_axi_awid[1]),
        .s1_axi_awaddr   (c0_axi_awaddr[1]),
        .s1_axi_awlen    (c0_axi_awlen[1]),
        .s1_axi_awsize   (c0_axi_awsize[1]),
        .s1_axi_awburst  (c0_axi_awburst[1]),
        .s1_axi_awlock   (c0_axi_awlock[1]),
        .s1_axi_awcache  (c0_axi_awcache[1]),
        .s1_axi_awprot   (c0_axi_awprot[1]),
        .s1_axi_awqos    (c0_axi_awqos[1]),
        .s1_axi_awvalid  (c0_axi_awvalid[1]),
        .s1_axi_awready  (c0_axi_awready[1]),
        .s1_axi_wdata    (c0_axi_wdata[1]),
        .s1_axi_wstrb    (c0_axi_wstrb[1]),
        .s1_axi_wlast    (c0_axi_wlast[1]),
        .s1_axi_wvalid   (c0_axi_wvalid[1]),
        .s1_axi_wready   (c0_axi_wready[1]),
        .s1_axi_bid      (c0_axi_bid[1]),
        .s1_axi_bresp    (c0_axi_bresp[1]),
        .s1_axi_bvalid   (c0_axi_bvalid[1]),
        .s1_axi_bready   (c0_axi_bready[1]),
        .s1_axi_arid     (c0_axi_arid[1]),
        .s1_axi_araddr   (c0_axi_araddr[1]),
        .s1_axi_arlen    (c0_axi_arlen[1]),
        .s1_axi_arsize   (c0_axi_arsize[1]),
        .s1_axi_arburst  (c0_axi_arburst[1]),
        .s1_axi_arlock   (c0_axi_arlock[1]),
        .s1_axi_arcache  (c0_axi_arcache[1]),
        .s1_axi_arprot   (c0_axi_arprot[1]),
        .s1_axi_arqos    (c0_axi_arqos[1]),
        .s1_axi_arvalid  (c0_axi_arvalid[1]),
        .s1_axi_arready  (c0_axi_arready[1]),
        .s1_axi_rid      (c0_axi_rid[1]),
        .s1_axi_rdata    (c0_axi_rdata[1]),
        .s1_axi_rresp    (c0_axi_rresp[1]),
        .s1_axi_rlast    (c0_axi_rlast[1]),
        .s1_axi_rvalid   (c0_axi_rvalid[1]),
        .s1_axi_rready   (c0_axi_rready[1]),
    `endif // PICO_AXI_PORT_1

   `ifdef PICO_AXI_PORT_2
        // master port 2
        .s2_axi_clk      (c0_axi_clk[2]),
        .s2_axi_awid     (c0_axi_awid[2]),
        .s2_axi_awaddr   (c0_axi_awaddr[2]),
        .s2_axi_awlen    (c0_axi_awlen[2]),
        .s2_axi_awsize   (c0_axi_awsize[2]),
        .s2_axi_awburst  (c0_axi_awburst[2]),
        .s2_axi_awlock   (c0_axi_awlock[2]),
        .s2_axi_awcache  (c0_axi_awcache[2]),
        .s2_axi_awprot   (c0_axi_awprot[2]),
        .s2_axi_awqos    (c0_axi_awqos[2]),
        .s2_axi_awvalid  (c0_axi_awvalid[2]),
        .s2_axi_awready  (c0_axi_awready[2]),
        .s2_axi_wdata    (c0_axi_wdata[2]),
        .s2_axi_wstrb    (c0_axi_wstrb[2]),
        .s2_axi_wlast    (c0_axi_wlast[2]),
        .s2_axi_wvalid   (c0_axi_wvalid[2]),
        .s2_axi_wready   (c0_axi_wready[2]),
        .s2_axi_bid      (c0_axi_bid[2]),
        .s2_axi_bresp    (c0_axi_bresp[2]),
        .s2_axi_bvalid   (c0_axi_bvalid[2]),
        .s2_axi_bready   (c0_axi_bready[2]),
        .s2_axi_arid     (c0_axi_arid[2]),
        .s2_axi_araddr   (c0_axi_araddr[2]),
        .s2_axi_arlen    (c0_axi_arlen[2]),
        .s2_axi_arsize   (c0_axi_arsize[2]),
        .s2_axi_arburst  (c0_axi_arburst[2]),
        .s2_axi_arlock   (c0_axi_arlock[2]),
        .s2_axi_arcache  (c0_axi_arcache[2]),
        .s2_axi_arprot   (c0_axi_arprot[2]),
        .s2_axi_arqos    (c0_axi_arqos[2]),
        .s2_axi_arvalid  (c0_axi_arvalid[2]),
        .s2_axi_arready  (c0_axi_arready[2]),
        .s2_axi_rid      (c0_axi_rid[2]),
        .s2_axi_rdata    (c0_axi_rdata[2]),
        .s2_axi_rresp    (c0_axi_rresp[2]),
        .s2_axi_rlast    (c0_axi_rlast[2]),
        .s2_axi_rvalid   (c0_axi_rvalid[2]),
        .s2_axi_rready   (c0_axi_rready[2]),
    `endif // PICO_AXI_PORT_2

   `ifdef PICO_AXI_PORT_3
        // master port 3
        .s3_axi_clk      (c0_axi_clk[3]),
        .s3_axi_awid     (c0_axi_awid[3]),
        .s3_axi_awaddr   (c0_axi_awaddr[3]),
        .s3_axi_awlen    (c0_axi_awlen[3]),
        .s3_axi_awsize   (c0_axi_awsize[3]),
        .s3_axi_awburst  (c0_axi_awburst[3]),
        .s3_axi_awlock   (c0_axi_awlock[3]),
        .s3_axi_awcache  (c0_axi_awcache[3]),
        .s3_axi_awprot   (c0_axi_awprot[3]),
        .s3_axi_awqos    (c0_axi_awqos[3]),
        .s3_axi_awvalid  (c0_axi_awvalid[3]),
        .s3_axi_awready  (c0_axi_awready[3]),
        .s3_axi_wdata    (c0_axi_wdata[3]),
        .s3_axi_wstrb    (c0_axi_wstrb[3]),
        .s3_axi_wlast    (c0_axi_wlast[3]),
        .s3_axi_wvalid   (c0_axi_wvalid[3]),
        .s3_axi_wready   (c0_axi_wready[3]),
        .s3_axi_bid      (c0_axi_bid[3]),
        .s3_axi_bresp    (c0_axi_bresp[3]),
        .s3_axi_bvalid   (c0_axi_bvalid[3]),
        .s3_axi_bready   (c0_axi_bready[3]),
        .s3_axi_arid     (c0_axi_arid[3]),
        .s3_axi_araddr   (c0_axi_araddr[3]),
        .s3_axi_arlen    (c0_axi_arlen[3]),
        .s3_axi_arsize   (c0_axi_arsize[3]),
        .s3_axi_arburst  (c0_axi_arburst[3]),
        .s3_axi_arlock   (c0_axi_arlock[3]),
        .s3_axi_arcache  (c0_axi_arcache[3]),
        .s3_axi_arprot   (c0_axi_arprot[3]),
        .s3_axi_arqos    (c0_axi_arqos[3]),
        .s3_axi_arvalid  (c0_axi_arvalid[3]),
        .s3_axi_arready  (c0_axi_arready[3]),
        .s3_axi_rid      (c0_axi_rid[3]),
        .s3_axi_rdata    (c0_axi_rdata[3]),
        .s3_axi_rresp    (c0_axi_rresp[3]),
        .s3_axi_rlast    (c0_axi_rlast[3]),
        .s3_axi_rvalid   (c0_axi_rvalid[3]),
        .s3_axi_rready   (c0_axi_rready[3]),
    `endif // PICO_AXI_PORT_3

   `ifdef PICO_AXI_PORT_4
        // master port 4
        .s4_axi_clk      (c0_axi_clk[4]),
        .s4_axi_awid     (c0_axi_awid[4]),
        .s4_axi_awaddr   (c0_axi_awaddr[4]),
        .s4_axi_awlen    (c0_axi_awlen[4]),
        .s4_axi_awsize   (c0_axi_awsize[4]),
        .s4_axi_awburst  (c0_axi_awburst[4]),
        .s4_axi_awlock   (c0_axi_awlock[4]),
        .s4_axi_awcache  (c0_axi_awcache[4]),
        .s4_axi_awprot   (c0_axi_awprot[4]),
        .s4_axi_awqos    (c0_axi_awqos[4]),
        .s4_axi_awvalid  (c0_axi_awvalid[4]),
        .s4_axi_awready  (c0_axi_awready[4]),
        .s4_axi_wdata    (c0_axi_wdata[4]),
        .s4_axi_wstrb    (c0_axi_wstrb[4]),
        .s4_axi_wlast    (c0_axi_wlast[4]),
        .s4_axi_wvalid   (c0_axi_wvalid[4]),
        .s4_axi_wready   (c0_axi_wready[4]),
        .s4_axi_bid      (c0_axi_bid[4]),
        .s4_axi_bresp    (c0_axi_bresp[4]),
        .s4_axi_bvalid   (c0_axi_bvalid[4]),
        .s4_axi_bready   (c0_axi_bready[4]),
        .s4_axi_arid     (c0_axi_arid[4]),
        .s4_axi_araddr   (c0_axi_araddr[4]),
        .s4_axi_arlen    (c0_axi_arlen[4]),
        .s4_axi_arsize   (c0_axi_arsize[4]),
        .s4_axi_arburst  (c0_axi_arburst[4]),
        .s4_axi_arlock   (c0_axi_arlock[4]),
        .s4_axi_arcache  (c0_axi_arcache[4]),
        .s4_axi_arprot   (c0_axi_arprot[4]),
        .s4_axi_arqos    (c0_axi_arqos[4]),
        .s4_axi_arvalid  (c0_axi_arvalid[4]),
        .s4_axi_arready  (c0_axi_arready[4]),
        .s4_axi_rid      (c0_axi_rid[4]),
        .s4_axi_rdata    (c0_axi_rdata[4]),
        .s4_axi_rresp    (c0_axi_rresp[4]),
        .s4_axi_rlast    (c0_axi_rlast[4]),
        .s4_axi_rvalid   (c0_axi_rvalid[4]),
        .s4_axi_rready   (c0_axi_rready[4]),
    `endif // PICO_AXI_PORT_4

   `ifdef PICO_AXI_PORT_5
        // master port 5
        .s5_axi_clk      (c0_axi_clk[5]),
        .s5_axi_awid     (c0_axi_awid[5]),
        .s5_axi_awaddr   (c0_axi_awaddr[5]),
        .s5_axi_awlen    (c0_axi_awlen[5]),
        .s5_axi_awsize   (c0_axi_awsize[5]),
        .s5_axi_awburst  (c0_axi_awburst[5]),
        .s5_axi_awlock   (c0_axi_awlock[5]),
        .s5_axi_awcache  (c0_axi_awcache[5]),
        .s5_axi_awprot   (c0_axi_awprot[5]),
        .s5_axi_awqos    (c0_axi_awqos[5]),
        .s5_axi_awvalid  (c0_axi_awvalid[5]),
        .s5_axi_awready  (c0_axi_awready[5]),
        .s5_axi_wdata    (c0_axi_wdata[5]),
        .s5_axi_wstrb    (c0_axi_wstrb[5]),
        .s5_axi_wlast    (c0_axi_wlast[5]),
        .s5_axi_wvalid   (c0_axi_wvalid[5]),
        .s5_axi_wready   (c0_axi_wready[5]),
        .s5_axi_bid      (c0_axi_bid[5]),
        .s5_axi_bresp    (c0_axi_bresp[5]),
        .s5_axi_bvalid   (c0_axi_bvalid[5]),
        .s5_axi_bready   (c0_axi_bready[5]),
        .s5_axi_arid     (c0_axi_arid[5]),
        .s5_axi_araddr   (c0_axi_araddr[5]),
        .s5_axi_arlen    (c0_axi_arlen[5]),
        .s5_axi_arsize   (c0_axi_arsize[5]),
        .s5_axi_arburst  (c0_axi_arburst[5]),
        .s5_axi_arlock   (c0_axi_arlock[5]),
        .s5_axi_arcache  (c0_axi_arcache[5]),
        .s5_axi_arprot   (c0_axi_arprot[5]),
        .s5_axi_arqos    (c0_axi_arqos[5]),
        .s5_axi_arvalid  (c0_axi_arvalid[5]),
        .s5_axi_arready  (c0_axi_arready[5]),
        .s5_axi_rid      (c0_axi_rid[5]),
        .s5_axi_rdata    (c0_axi_rdata[5]),
        .s5_axi_rresp    (c0_axi_rresp[5]),
        .s5_axi_rlast    (c0_axi_rlast[5]),
        .s5_axi_rvalid   (c0_axi_rvalid[5]),
        .s5_axi_rready   (c0_axi_rready[5]),
    `endif // PICO_AXI_PORT_5

   `ifdef PICO_AXI_PORT_6
        // master port 6
        .s6_axi_clk      (c0_axi_clk[6]),
        .s6_axi_awid     (c0_axi_awid[6]),
        .s6_axi_awaddr   (c0_axi_awaddr[6]),
        .s6_axi_awlen    (c0_axi_awlen[6]),
        .s6_axi_awsize   (c0_axi_awsize[6]),
        .s6_axi_awburst  (c0_axi_awburst[6]),
        .s6_axi_awlock   (c0_axi_awlock[6]),
        .s6_axi_awcache  (c0_axi_awcache[6]),
        .s6_axi_awprot   (c0_axi_awprot[6]),
        .s6_axi_awqos    (c0_axi_awqos[6]),
        .s6_axi_awvalid  (c0_axi_awvalid[6]),
        .s6_axi_awready  (c0_axi_awready[6]),
        .s6_axi_wdata    (c0_axi_wdata[6]),
        .s6_axi_wstrb    (c0_axi_wstrb[6]),
        .s6_axi_wlast    (c0_axi_wlast[6]),
        .s6_axi_wvalid   (c0_axi_wvalid[6]),
        .s6_axi_wready   (c0_axi_wready[6]),
        .s6_axi_bid      (c0_axi_bid[6]),
        .s6_axi_bresp    (c0_axi_bresp[6]),
        .s6_axi_bvalid   (c0_axi_bvalid[6]),
        .s6_axi_bready   (c0_axi_bready[6]),
        .s6_axi_arid     (c0_axi_arid[6]),
        .s6_axi_araddr   (c0_axi_araddr[6]),
        .s6_axi_arlen    (c0_axi_arlen[6]),
        .s6_axi_arsize   (c0_axi_arsize[6]),
        .s6_axi_arburst  (c0_axi_arburst[6]),
        .s6_axi_arlock   (c0_axi_arlock[6]),
        .s6_axi_arcache  (c0_axi_arcache[6]),
        .s6_axi_arprot   (c0_axi_arprot[6]),
        .s6_axi_arqos    (c0_axi_arqos[6]),
        .s6_axi_arvalid  (c0_axi_arvalid[6]),
        .s6_axi_arready  (c0_axi_arready[6]),
        .s6_axi_rid      (c0_axi_rid[6]),
        .s6_axi_rdata    (c0_axi_rdata[6]),
        .s6_axi_rresp    (c0_axi_rresp[6]),
        .s6_axi_rlast    (c0_axi_rlast[6]),
        .s6_axi_rvalid   (c0_axi_rvalid[6]),
        .s6_axi_rready   (c0_axi_rready[6]),
    `endif // PICO_AXI_PORT_6

   `ifdef PICO_AXI_PORT_7
        // master port 7
        .s7_axi_clk      (c0_axi_clk[7]),
        .s7_axi_awid     (c0_axi_awid[7]),
        .s7_axi_awaddr   (c0_axi_awaddr[7]),
        .s7_axi_awlen    (c0_axi_awlen[7]),
        .s7_axi_awsize   (c0_axi_awsize[7]),
        .s7_axi_awburst  (c0_axi_awburst[7]),
        .s7_axi_awlock   (c0_axi_awlock[7]),
        .s7_axi_awcache  (c0_axi_awcache[7]),
        .s7_axi_awprot   (c0_axi_awprot[7]),
        .s7_axi_awqos    (c0_axi_awqos[7]),
        .s7_axi_awvalid  (c0_axi_awvalid[7]),
        .s7_axi_awready  (c0_axi_awready[7]),
        .s7_axi_wdata    (c0_axi_wdata[7]),
        .s7_axi_wstrb    (c0_axi_wstrb[7]),
        .s7_axi_wlast    (c0_axi_wlast[7]),
        .s7_axi_wvalid   (c0_axi_wvalid[7]),
        .s7_axi_wready   (c0_axi_wready[7]),
        .s7_axi_bid      (c0_axi_bid[7]),
        .s7_axi_bresp    (c0_axi_bresp[7]),
        .s7_axi_bvalid   (c0_axi_bvalid[7]),
        .s7_axi_bready   (c0_axi_bready[7]),
        .s7_axi_arid     (c0_axi_arid[7]),
        .s7_axi_araddr   (c0_axi_araddr[7]),
        .s7_axi_arlen    (c0_axi_arlen[7]),
        .s7_axi_arsize   (c0_axi_arsize[7]),
        .s7_axi_arburst  (c0_axi_arburst[7]),
        .s7_axi_arlock   (c0_axi_arlock[7]),
        .s7_axi_arcache  (c0_axi_arcache[7]),
        .s7_axi_arprot   (c0_axi_arprot[7]),
        .s7_axi_arqos    (c0_axi_arqos[7]),
        .s7_axi_arvalid  (c0_axi_arvalid[7]),
        .s7_axi_arready  (c0_axi_arready[7]),
        .s7_axi_rid      (c0_axi_rid[7]),
        .s7_axi_rdata    (c0_axi_rdata[7]),
        .s7_axi_rresp    (c0_axi_rresp[7]),
        .s7_axi_rlast    (c0_axi_rlast[7]),
        .s7_axi_rvalid   (c0_axi_rvalid[7]),
        .s7_axi_rready   (c0_axi_rready[7]),
    `endif // PICO_AXI_PORT_7


    `ifdef ALTERA_FPGA
        //avalon interface
        .avl_ready         (avl_ready),
        .avl_addr          (avl_addr),
        .avl_rdata_valid   (avl_rdata_valid),
        .avl_rdata         (avl_rdata),
        .avl_wdata         (avl_wdata),
        .avl_be            (avl_be),
        .avl_read_req      (avl_read_req),
        .avl_write_req     (avl_write_req),
        .avl_size          (avl_size)
    `else
        .m_axi_awid         (c0_s_axi_awid),
        .m_axi_awaddr       (c0_s_axi_awaddr),
        .m_axi_awlen        (c0_s_axi_awlen),
        .m_axi_awsize       (c0_s_axi_awsize),
        .m_axi_awburst      (c0_s_axi_awburst),
        .m_axi_awlock       (c0_s_axi_awlock),
        .m_axi_awcache      (c0_s_axi_awcache),
        .m_axi_awprot       (c0_s_axi_awprot),
        .m_axi_awqos        (c0_s_axi_awqos),
        .m_axi_awvalid      (c0_s_axi_awvalid),
        .m_axi_awready      (c0_s_axi_awready),
        .m_axi_wdata        (c0_s_axi_wdata),
        .m_axi_wstrb        (c0_s_axi_wstrb),
        .m_axi_wlast        (c0_s_axi_wlast),
        .m_axi_wvalid       (c0_s_axi_wvalid),
        .m_axi_wready       (c0_s_axi_wready),
        .m_axi_bid          (c0_s_axi_bid),
        .m_axi_bresp        (c0_s_axi_bresp),
        .m_axi_bvalid       (c0_s_axi_bvalid),
        .m_axi_bready       (c0_s_axi_bready),
        .m_axi_arid         (c0_s_axi_arid),
        .m_axi_araddr       (c0_s_axi_araddr),
        .m_axi_arlen        (c0_s_axi_arlen),
        .m_axi_arsize       (c0_s_axi_arsize),
        .m_axi_arburst      (c0_s_axi_arburst),
        .m_axi_arlock       (c0_s_axi_arlock),
        .m_axi_arcache      (c0_s_axi_arcache),
        .m_axi_arprot       (c0_s_axi_arprot),
        .m_axi_arqos        (c0_s_axi_arqos),
        .m_axi_arvalid      (c0_s_axi_arvalid),
        .m_axi_arready      (c0_s_axi_arready),
        .m_axi_rid          (c0_s_axi_rid),
        .m_axi_rdata        (c0_s_axi_rdata),
        .m_axi_rresp        (c0_s_axi_rresp),
        .m_axi_rlast        (c0_s_axi_rlast),
        .m_axi_rvalid       (c0_s_axi_rvalid),
        .m_axi_rready       (c0_s_axi_rready)
    `endif // ALTERA_FPGA
    );

    assign c0_axi_clk[0] = clk;
`endif


    /////////////////////////
    // Stream Controller 0 //
    /////////////////////////
    // host streaming interface sits on port 0 of the axi interconnect
    PicoStreamToAXI #(
        .C_AXI_ID_WIDTH     (C0_C_S_AXI_ID_WIDTH-4),
        .C_AXI_ADDR_WIDTH   (C0_C_S_AXI_ADDR_WIDTH),
        .STREAM_DATA_WIDTH  (128),
        .UPSIZE_RATIO       (C0_C_S_AXI_DATA_WIDTH/128),
        .LOG_UPSIZE_RATIO   (clogb2(C0_C_S_AXI_DATA_WIDTH/128))
    )
    stream_to_mem_0
    (
        // streaming interface
        .clk                (clk),
        .rst                (rst),

`ifdef PICO_DDR3
        .si_ready           (stream_in_rdy[`DDR3_STREAM_ID]),
        .si_valid           (stream_in_valid[`DDR3_STREAM_ID]),
        .si_data            (stream_in_data[`DDR3_STREAM_ID][127:0]),
        .so_ready           (stream_out_rdy[`DDR3_STREAM_ID]),
        .so_valid           (stream_out_valid[`DDR3_STREAM_ID]),
        .so_data            (stream_out_data[`DDR3_STREAM_ID][127:0]),
`elsif PICO_DDR4
        .si_ready           (stream_in_rdy[`DDR4_STREAM_ID]),
        .si_valid           (stream_in_valid[`DDR4_STREAM_ID]),
        .si_data            (stream_in_data[`DDR4_STREAM_ID][127:0]),
        .so_ready           (stream_out_rdy[`DDR4_STREAM_ID]),
        .so_valid           (stream_out_valid[`DDR4_STREAM_ID]),
        .so_data            (stream_out_data[`DDR4_STREAM_ID][127:0]),
`endif // PICO_DDR

        // ddr3 signals
        .ddr3_reset         (ddr3_sys_rst[0]),
        .init_cmptd         (c0_phy_init_done),

        // axi interface
        .s_axi_awid         (c0_axi_awid[0]),
        .s_axi_awaddr       (c0_axi_awaddr[0]),
        .s_axi_awlen        (c0_axi_awlen[0]),
        .s_axi_awsize       (c0_axi_awsize[0]),
        .s_axi_awburst      (c0_axi_awburst[0]),
        .s_axi_awlock       (c0_axi_awlock[0]),
        .s_axi_awcache      (c0_axi_awcache[0]),
        .s_axi_awprot       (c0_axi_awprot[0]),
        .s_axi_awqos        (c0_axi_awqos[0]),
        .s_axi_awvalid      (c0_axi_awvalid[0]),
        .s_axi_awready      (c0_axi_awready[0]),
        .s_axi_wdata        (c0_axi_wdata[0]),
        .s_axi_wstrb        (c0_axi_wstrb[0]),
        .s_axi_wlast        (c0_axi_wlast[0]),
        .s_axi_wvalid       (c0_axi_wvalid[0]),
        .s_axi_wready       (c0_axi_wready[0]),
        .s_axi_bid          (c0_axi_bid[0]),
        .s_axi_bresp        (c0_axi_bresp[0]),
        .s_axi_bvalid       (c0_axi_bvalid[0]),
        .s_axi_bready       (c0_axi_bready[0]),
        .s_axi_arid         (c0_axi_arid[0]),
        .s_axi_araddr       (c0_axi_araddr[0]),
        .s_axi_arlen        (c0_axi_arlen[0]),
        .s_axi_arsize       (c0_axi_arsize[0]),
        .s_axi_arburst      (c0_axi_arburst[0]),
        .s_axi_arlock       (c0_axi_arlock[0]),
        .s_axi_arcache      (c0_axi_arcache[0]),
        .s_axi_arprot       (c0_axi_arprot[0]),
        .s_axi_arqos        (c0_axi_arqos[0]),
        .s_axi_arvalid      (c0_axi_arvalid[0]),
        .s_axi_arready      (c0_axi_arready[0]),
        .s_axi_rid          (c0_axi_rid[0]),
        .s_axi_rdata        (c0_axi_rdata[0]),
        .s_axi_rresp        (c0_axi_rresp[0]),
        .s_axi_rlast        (c0_axi_rlast[0]),
        .s_axi_rvalid       (c0_axi_rvalid[0]),
        .s_axi_rready       (c0_axi_rready[0])
    );

`endif// PICO_DDR3_OR_DDR4

    `ifdef PICOBUS_WIDTH                 // Only enable these streams if there is a User module using the picobus

        Stream2PicoBus #(
	    .STREAM_ID(125),
	    .W(`PICOBUS_WIDTH),
	    .C_DATA_WIDTH(C_DATA_WIDTH),
	    .S_PB_RATIO(S_PB_RATIO)
        ) UserModule_s2pb (
            .s_clk(clk),
            .s_rst(rst),

            .s_out_en(s_out_en),
            .s_out_id(s_out_id),
            .s_out_data(s_out_data_userpb),
	    .s_out_ow_dvld(s_out_ow_dvld_userpb),

            .s_in_valid(s_in_valid),
            .s_in_id(s_in_id[8:0]),
            .s_in_data(s_in_data[C_DATA_WIDTH-1:0]),
	    .s_in_ow_dvld(s_in_ow_dvld[OW_DVLD_W-1:0]),

            .s_poll_id(s_poll_id[8:0]),
            .s_poll_seq(s_poll_seq_userpb[31:0]),
            .s_poll_next_desc(s_poll_next_desc_userpb[127:0]),
            .s_poll_next_desc_valid(s_poll_next_desc_valid_userpb),

            .s_next_desc_rd_en(s_next_desc_rd_en),
            .s_next_desc_rd_id(s_next_desc_rd_id[8:0]),

            .PicoClk(UserModulePicoClk),
            .PicoRst(UserModulePicoRst),
            .PicoWr(UserModulePicoWr),
            .PicoDataIn(UserModulePicoDataIn),
            .PicoRd(UserModulePicoRd),
            .PicoAddr(UserModulePicoAddr),
            .PicoDataOut(UserModulePicoDataOut `ifdef ENABLE_HMC | PicoDataOut `endif)
        );
    `endif // PICOBUS_WIDTH

    // begin usermodule Stream Interface

    localparam INSTREAM = {72'h0
                `ifdef STREAM1_IN_WIDTH `ifdef STREAM1_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM1_IN_WIDTH , 8'd1 `endif
                `ifdef STREAM2_IN_WIDTH `ifdef STREAM2_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM2_IN_WIDTH , 8'd2 `endif
                `ifdef STREAM3_IN_WIDTH `ifdef STREAM3_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM3_IN_WIDTH , 8'd3 `endif
                `ifdef STREAM4_IN_WIDTH `ifdef STREAM4_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM4_IN_WIDTH , 8'd4 `endif
                `ifdef STREAM5_IN_WIDTH `ifdef STREAM5_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM5_IN_WIDTH , 8'd5 `endif
                `ifdef STREAM6_IN_WIDTH `ifdef STREAM6_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM6_IN_WIDTH , 8'd6 `endif
                `ifdef STREAM7_IN_WIDTH `ifdef STREAM7_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM7_IN_WIDTH , 8'd7 `endif
                `ifdef STREAM8_IN_WIDTH `ifdef STREAM8_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM8_IN_WIDTH , 8'd8 `endif
                `ifdef STREAM9_IN_WIDTH `ifdef STREAM9_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM9_IN_WIDTH , 8'd9 `endif
                `ifdef STREAM10_IN_WIDTH `ifdef STREAM10_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM10_IN_WIDTH , 8'd10 `endif
                `ifdef STREAM11_IN_WIDTH `ifdef STREAM11_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM11_IN_WIDTH , 8'd11 `endif
                `ifdef STREAM12_IN_WIDTH `ifdef STREAM12_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM12_IN_WIDTH , 8'd12 `endif
                `ifdef STREAM13_IN_WIDTH `ifdef STREAM13_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM13_IN_WIDTH , 8'd13 `endif
                `ifdef STREAM14_IN_WIDTH `ifdef STREAM14_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM14_IN_WIDTH , 8'd14 `endif
                `ifdef STREAM15_IN_WIDTH `ifdef STREAM15_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM15_IN_WIDTH , 8'd15 `endif
                `ifdef STREAM16_IN_WIDTH `ifdef STREAM16_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM16_IN_WIDTH , 8'd16 `endif
                `ifdef STREAM17_IN_WIDTH `ifdef STREAM17_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM17_IN_WIDTH , 8'd17 `endif
                `ifdef STREAM18_IN_WIDTH `ifdef STREAM18_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM18_IN_WIDTH , 8'd18 `endif
                `ifdef STREAM19_IN_WIDTH `ifdef STREAM19_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM19_IN_WIDTH , 8'd19 `endif
                `ifdef STREAM20_IN_WIDTH `ifdef STREAM20_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM20_IN_WIDTH , 8'd20 `endif
                `ifdef STREAM21_IN_WIDTH `ifdef STREAM21_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM21_IN_WIDTH , 8'd21 `endif
                `ifdef STREAM22_IN_WIDTH `ifdef STREAM22_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM22_IN_WIDTH , 8'd22 `endif
                `ifdef STREAM23_IN_WIDTH `ifdef STREAM23_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM23_IN_WIDTH , 8'd23 `endif
                `ifdef STREAM24_IN_WIDTH `ifdef STREAM24_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM24_IN_WIDTH , 8'd24 `endif
                `ifdef STREAM25_IN_WIDTH `ifdef STREAM25_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM25_IN_WIDTH , 8'd25 `endif
                `ifdef STREAM26_IN_WIDTH `ifdef STREAM26_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM26_IN_WIDTH , 8'd26 `endif
                `ifdef STREAM27_IN_WIDTH `ifdef STREAM27_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM27_IN_WIDTH , 8'd27 `endif
                `ifdef STREAM28_IN_WIDTH `ifdef STREAM28_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM28_IN_WIDTH , 8'd28 `endif
                `ifdef STREAM29_IN_WIDTH `ifdef STREAM29_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM29_IN_WIDTH , 8'd29 `endif
                `ifdef STREAM30_IN_WIDTH `ifdef STREAM30_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM30_IN_WIDTH , 8'd30 `endif
                `ifdef STREAM31_IN_WIDTH `ifdef STREAM31_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM31_IN_WIDTH , 8'd31 `endif
                `ifdef STREAM32_IN_WIDTH `ifdef STREAM32_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM32_IN_WIDTH , 8'd32 `endif
                `ifdef STREAM33_IN_WIDTH `ifdef STREAM33_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM33_IN_WIDTH , 8'd33 `endif
                `ifdef STREAM34_IN_WIDTH `ifdef STREAM34_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM34_IN_WIDTH , 8'd34 `endif
                `ifdef STREAM35_IN_WIDTH `ifdef STREAM35_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM35_IN_WIDTH , 8'd35 `endif
                `ifdef STREAM36_IN_WIDTH `ifdef STREAM36_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM36_IN_WIDTH , 8'd36 `endif
                `ifdef STREAM37_IN_WIDTH `ifdef STREAM37_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM37_IN_WIDTH , 8'd37 `endif
                `ifdef STREAM38_IN_WIDTH `ifdef STREAM38_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM38_IN_WIDTH , 8'd38 `endif
                `ifdef STREAM39_IN_WIDTH `ifdef STREAM39_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM39_IN_WIDTH , 8'd39 `endif
                `ifdef STREAM40_IN_WIDTH `ifdef STREAM40_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM40_IN_WIDTH , 8'd40 `endif
                `ifdef STREAM41_IN_WIDTH `ifdef STREAM41_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM41_IN_WIDTH , 8'd41 `endif
                `ifdef STREAM42_IN_WIDTH `ifdef STREAM42_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM42_IN_WIDTH , 8'd42 `endif
                `ifdef STREAM43_IN_WIDTH `ifdef STREAM43_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM43_IN_WIDTH , 8'd43 `endif
                `ifdef STREAM44_IN_WIDTH `ifdef STREAM44_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM44_IN_WIDTH , 8'd44 `endif
                `ifdef STREAM45_IN_WIDTH `ifdef STREAM45_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM45_IN_WIDTH , 8'd45 `endif
                `ifdef STREAM46_IN_WIDTH `ifdef STREAM46_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM46_IN_WIDTH , 8'd46 `endif
                `ifdef STREAM47_IN_WIDTH `ifdef STREAM47_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM47_IN_WIDTH , 8'd47 `endif
                `ifdef STREAM48_IN_WIDTH `ifdef STREAM48_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM48_IN_WIDTH , 8'd48 `endif
                `ifdef STREAM49_IN_WIDTH `ifdef STREAM49_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM49_IN_WIDTH , 8'd49 `endif
                `ifdef STREAM50_IN_WIDTH `ifdef STREAM50_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM50_IN_WIDTH , 8'd50 `endif
                `ifdef STREAM51_IN_WIDTH `ifdef STREAM51_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM51_IN_WIDTH , 8'd51 `endif
                `ifdef STREAM52_IN_WIDTH `ifdef STREAM52_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM52_IN_WIDTH , 8'd52 `endif
                `ifdef STREAM53_IN_WIDTH `ifdef STREAM53_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM53_IN_WIDTH , 8'd53 `endif
                `ifdef STREAM54_IN_WIDTH `ifdef STREAM54_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM54_IN_WIDTH , 8'd54 `endif
                `ifdef STREAM55_IN_WIDTH `ifdef STREAM55_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM55_IN_WIDTH , 8'd55 `endif
                `ifdef STREAM56_IN_WIDTH `ifdef STREAM56_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM56_IN_WIDTH , 8'd56 `endif
                `ifdef STREAM57_IN_WIDTH `ifdef STREAM57_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM57_IN_WIDTH , 8'd57 `endif
                `ifdef STREAM58_IN_WIDTH `ifdef STREAM58_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM58_IN_WIDTH , 8'd58 `endif
                `ifdef STREAM59_IN_WIDTH `ifdef STREAM59_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM59_IN_WIDTH , 8'd59 `endif
                `ifdef STREAM60_IN_WIDTH `ifdef STREAM60_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM60_IN_WIDTH , 8'd60 `endif
                `ifdef STREAM61_IN_WIDTH `ifdef STREAM61_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM61_IN_WIDTH , 8'd61 `endif
                `ifdef STREAM62_IN_WIDTH `ifdef STREAM62_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM62_IN_WIDTH , 8'd62 `endif
                `ifdef STREAM63_IN_WIDTH `ifdef STREAM63_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM63_IN_WIDTH , 8'd63 `endif
                `ifdef STREAM64_IN_WIDTH `ifdef STREAM64_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM64_IN_WIDTH , 8'd64 `endif
                `ifdef STREAM65_IN_WIDTH `ifdef STREAM65_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM65_IN_WIDTH , 8'd65 `endif
                `ifdef STREAM66_IN_WIDTH `ifdef STREAM66_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM66_IN_WIDTH , 8'd66 `endif
                `ifdef STREAM67_IN_WIDTH `ifdef STREAM67_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM67_IN_WIDTH , 8'd67 `endif
                `ifdef STREAM68_IN_WIDTH `ifdef STREAM68_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM68_IN_WIDTH , 8'd68 `endif
                `ifdef STREAM69_IN_WIDTH `ifdef STREAM69_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM69_IN_WIDTH , 8'd69 `endif
                `ifdef STREAM70_IN_WIDTH `ifdef STREAM70_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM70_IN_WIDTH , 8'd70 `endif
                `ifdef STREAM71_IN_WIDTH `ifdef STREAM71_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM71_IN_WIDTH , 8'd71 `endif
                `ifdef STREAM72_IN_WIDTH `ifdef STREAM72_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM72_IN_WIDTH , 8'd72 `endif
                `ifdef STREAM73_IN_WIDTH `ifdef STREAM73_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM73_IN_WIDTH , 8'd73 `endif
                `ifdef STREAM74_IN_WIDTH `ifdef STREAM74_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM74_IN_WIDTH , 8'd74 `endif
                `ifdef STREAM75_IN_WIDTH `ifdef STREAM75_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM75_IN_WIDTH , 8'd75 `endif
                `ifdef STREAM76_IN_WIDTH `ifdef STREAM76_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM76_IN_WIDTH , 8'd76 `endif
                `ifdef STREAM77_IN_WIDTH `ifdef STREAM77_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM77_IN_WIDTH , 8'd77 `endif
                `ifdef STREAM78_IN_WIDTH `ifdef STREAM78_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM78_IN_WIDTH , 8'd78 `endif
                `ifdef STREAM79_IN_WIDTH `ifdef STREAM79_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM79_IN_WIDTH , 8'd79 `endif
                `ifdef STREAM80_IN_WIDTH `ifdef STREAM80_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM80_IN_WIDTH , 8'd80 `endif
                `ifdef STREAM81_IN_WIDTH `ifdef STREAM81_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM81_IN_WIDTH , 8'd81 `endif
                `ifdef STREAM82_IN_WIDTH `ifdef STREAM82_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM82_IN_WIDTH , 8'd82 `endif
                `ifdef STREAM83_IN_WIDTH `ifdef STREAM83_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM83_IN_WIDTH , 8'd83 `endif
                `ifdef STREAM84_IN_WIDTH `ifdef STREAM84_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM84_IN_WIDTH , 8'd84 `endif
                `ifdef STREAM85_IN_WIDTH `ifdef STREAM85_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM85_IN_WIDTH , 8'd85 `endif
                `ifdef STREAM86_IN_WIDTH `ifdef STREAM86_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM86_IN_WIDTH , 8'd86 `endif
                `ifdef STREAM87_IN_WIDTH `ifdef STREAM87_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM87_IN_WIDTH , 8'd87 `endif
                `ifdef STREAM88_IN_WIDTH `ifdef STREAM88_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM88_IN_WIDTH , 8'd88 `endif
                `ifdef STREAM89_IN_WIDTH `ifdef STREAM89_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM89_IN_WIDTH , 8'd89 `endif
                `ifdef STREAM90_IN_WIDTH `ifdef STREAM90_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM90_IN_WIDTH , 8'd90 `endif
                `ifdef STREAM91_IN_WIDTH `ifdef STREAM91_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM91_IN_WIDTH , 8'd91 `endif
                `ifdef STREAM92_IN_WIDTH `ifdef STREAM92_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM92_IN_WIDTH , 8'd92 `endif
                `ifdef STREAM93_IN_WIDTH `ifdef STREAM93_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM93_IN_WIDTH , 8'd93 `endif
                `ifdef STREAM94_IN_WIDTH `ifdef STREAM94_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM94_IN_WIDTH , 8'd94 `endif
                `ifdef STREAM95_IN_WIDTH `ifdef STREAM95_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM95_IN_WIDTH , 8'd95 `endif
                `ifdef STREAM96_IN_WIDTH `ifdef STREAM96_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM96_IN_WIDTH , 8'd96 `endif
                `ifdef STREAM97_IN_WIDTH `ifdef STREAM97_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM97_IN_WIDTH , 8'd97 `endif
                `ifdef STREAM98_IN_WIDTH `ifdef STREAM98_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM98_IN_WIDTH , 8'd98 `endif
                `ifdef STREAM99_IN_WIDTH `ifdef STREAM99_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM99_IN_WIDTH , 8'd99 `endif
                `ifdef STREAM100_IN_WIDTH `ifdef STREAM100_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM100_IN_WIDTH , 8'd100 `endif
                `ifdef STREAM101_IN_WIDTH `ifdef STREAM101_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM101_IN_WIDTH , 8'd101 `endif
                `ifdef STREAM102_IN_WIDTH `ifdef STREAM102_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM102_IN_WIDTH , 8'd102 `endif
                `ifdef STREAM103_IN_WIDTH `ifdef STREAM103_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM103_IN_WIDTH , 8'd103 `endif
                `ifdef STREAM104_IN_WIDTH `ifdef STREAM104_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM104_IN_WIDTH , 8'd104 `endif
                `ifdef STREAM105_IN_WIDTH `ifdef STREAM105_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM105_IN_WIDTH , 8'd105 `endif
                `ifdef STREAM106_IN_WIDTH `ifdef STREAM106_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM106_IN_WIDTH , 8'd106 `endif
                `ifdef STREAM107_IN_WIDTH `ifdef STREAM107_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM107_IN_WIDTH , 8'd107 `endif
                `ifdef STREAM108_IN_WIDTH `ifdef STREAM108_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM108_IN_WIDTH , 8'd108 `endif
                `ifdef STREAM109_IN_WIDTH `ifdef STREAM109_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM109_IN_WIDTH , 8'd109 `endif
                `ifdef STREAM110_IN_WIDTH `ifdef STREAM110_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM110_IN_WIDTH , 8'd110 `endif
                `ifdef STREAM111_IN_WIDTH `ifdef STREAM111_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM111_IN_WIDTH , 8'd111 `endif
                `ifdef STREAM112_IN_WIDTH `ifdef STREAM112_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM112_IN_WIDTH , 8'd112 `endif
                `ifdef STREAM113_IN_WIDTH `ifdef STREAM113_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM113_IN_WIDTH , 8'd113 `endif
                `ifdef STREAM114_IN_WIDTH `ifdef STREAM114_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM114_IN_WIDTH , 8'd114 `endif
                `ifdef STREAM115_IN_WIDTH `ifdef STREAM115_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM115_IN_WIDTH , 8'd115 `endif
                `ifdef STREAM116_IN_WIDTH `ifdef STREAM116_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM116_IN_WIDTH , 8'd116 `endif
                `ifdef STREAM117_IN_WIDTH `ifdef STREAM117_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM117_IN_WIDTH , 8'd117 `endif
                `ifdef STREAM118_IN_WIDTH `ifdef STREAM118_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM118_IN_WIDTH , 8'd118 `endif
                `ifdef STREAM119_IN_WIDTH `ifdef STREAM119_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM119_IN_WIDTH , 8'd119 `endif
                `ifdef STREAM120_IN_WIDTH `ifdef STREAM120_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM120_IN_WIDTH , 8'd120 `endif
                `ifdef STREAM121_IN_WIDTH `ifdef STREAM121_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM121_IN_WIDTH , 8'd121 `endif
                `ifdef STREAM122_IN_WIDTH `ifdef STREAM122_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM122_IN_WIDTH , 8'd122 `endif
                `ifdef STREAM123_IN_WIDTH `ifdef STREAM123_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM123_IN_WIDTH , 8'd123 `endif
                `ifdef STREAM124_IN_WIDTH `ifdef STREAM124_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM124_IN_WIDTH , 8'd124 `endif
                `ifdef STREAM125_IN_WIDTH `ifdef STREAM125_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM125_IN_WIDTH , 8'd125 `endif
                `ifdef STREAM126_IN_WIDTH `ifdef STREAM126_IN_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM126_IN_WIDTH , 8'd126 `endif
                    };

    localparam OUTSTREAM = {72'h0
                `ifdef STREAM1_OUT_WIDTH `ifdef STREAM1_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM1_OUT_WIDTH , 8'd1 `endif
                `ifdef STREAM2_OUT_WIDTH `ifdef STREAM2_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM2_OUT_WIDTH , 8'd2 `endif
                `ifdef STREAM3_OUT_WIDTH `ifdef STREAM3_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM3_OUT_WIDTH , 8'd3 `endif
                `ifdef STREAM4_OUT_WIDTH `ifdef STREAM4_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM4_OUT_WIDTH , 8'd4 `endif
                `ifdef STREAM5_OUT_WIDTH `ifdef STREAM5_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM5_OUT_WIDTH , 8'd5 `endif
                `ifdef STREAM6_OUT_WIDTH `ifdef STREAM6_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM6_OUT_WIDTH , 8'd6 `endif
                `ifdef STREAM7_OUT_WIDTH `ifdef STREAM7_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM7_OUT_WIDTH , 8'd7 `endif
                `ifdef STREAM8_OUT_WIDTH `ifdef STREAM8_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM8_OUT_WIDTH , 8'd8 `endif
                `ifdef STREAM9_OUT_WIDTH `ifdef STREAM9_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM9_OUT_WIDTH , 8'd9 `endif
                `ifdef STREAM10_OUT_WIDTH `ifdef STREAM10_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM10_OUT_WIDTH , 8'd10 `endif
                `ifdef STREAM11_OUT_WIDTH `ifdef STREAM11_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM11_OUT_WIDTH , 8'd11 `endif
                `ifdef STREAM12_OUT_WIDTH `ifdef STREAM12_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM12_OUT_WIDTH , 8'd12 `endif
                `ifdef STREAM13_OUT_WIDTH `ifdef STREAM13_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM13_OUT_WIDTH , 8'd13 `endif
                `ifdef STREAM14_OUT_WIDTH `ifdef STREAM14_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM14_OUT_WIDTH , 8'd14 `endif
                `ifdef STREAM15_OUT_WIDTH `ifdef STREAM15_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM15_OUT_WIDTH , 8'd15 `endif
                `ifdef STREAM16_OUT_WIDTH `ifdef STREAM16_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM16_OUT_WIDTH , 8'd16 `endif
                `ifdef STREAM17_OUT_WIDTH `ifdef STREAM17_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM17_OUT_WIDTH , 8'd17 `endif
                `ifdef STREAM18_OUT_WIDTH `ifdef STREAM18_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM18_OUT_WIDTH , 8'd18 `endif
                `ifdef STREAM19_OUT_WIDTH `ifdef STREAM19_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM19_OUT_WIDTH , 8'd19 `endif
                `ifdef STREAM20_OUT_WIDTH `ifdef STREAM20_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM20_OUT_WIDTH , 8'd20 `endif
                `ifdef STREAM21_OUT_WIDTH `ifdef STREAM21_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM21_OUT_WIDTH , 8'd21 `endif
                `ifdef STREAM22_OUT_WIDTH `ifdef STREAM22_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM22_OUT_WIDTH , 8'd22 `endif
                `ifdef STREAM23_OUT_WIDTH `ifdef STREAM23_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM23_OUT_WIDTH , 8'd23 `endif
                `ifdef STREAM24_OUT_WIDTH `ifdef STREAM24_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM24_OUT_WIDTH , 8'd24 `endif
                `ifdef STREAM25_OUT_WIDTH `ifdef STREAM25_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM25_OUT_WIDTH , 8'd25 `endif
                `ifdef STREAM26_OUT_WIDTH `ifdef STREAM26_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM26_OUT_WIDTH , 8'd26 `endif
                `ifdef STREAM27_OUT_WIDTH `ifdef STREAM27_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM27_OUT_WIDTH , 8'd27 `endif
                `ifdef STREAM28_OUT_WIDTH `ifdef STREAM28_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM28_OUT_WIDTH , 8'd28 `endif
                `ifdef STREAM29_OUT_WIDTH `ifdef STREAM29_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM29_OUT_WIDTH , 8'd29 `endif
                `ifdef STREAM30_OUT_WIDTH `ifdef STREAM30_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM30_OUT_WIDTH , 8'd30 `endif
                `ifdef STREAM31_OUT_WIDTH `ifdef STREAM31_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM31_OUT_WIDTH , 8'd31 `endif
                `ifdef STREAM32_OUT_WIDTH `ifdef STREAM32_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM32_OUT_WIDTH , 8'd32 `endif
                `ifdef STREAM33_OUT_WIDTH `ifdef STREAM33_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM33_OUT_WIDTH , 8'd33 `endif
                `ifdef STREAM34_OUT_WIDTH `ifdef STREAM34_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM34_OUT_WIDTH , 8'd34 `endif
                `ifdef STREAM35_OUT_WIDTH `ifdef STREAM35_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM35_OUT_WIDTH , 8'd35 `endif
                `ifdef STREAM36_OUT_WIDTH `ifdef STREAM36_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM36_OUT_WIDTH , 8'd36 `endif
                `ifdef STREAM37_OUT_WIDTH `ifdef STREAM37_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM37_OUT_WIDTH , 8'd37 `endif
                `ifdef STREAM38_OUT_WIDTH `ifdef STREAM38_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM38_OUT_WIDTH , 8'd38 `endif
                `ifdef STREAM39_OUT_WIDTH `ifdef STREAM39_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM39_OUT_WIDTH , 8'd39 `endif
                `ifdef STREAM40_OUT_WIDTH `ifdef STREAM40_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM40_OUT_WIDTH , 8'd40 `endif
                `ifdef STREAM41_OUT_WIDTH `ifdef STREAM41_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM41_OUT_WIDTH , 8'd41 `endif
                `ifdef STREAM42_OUT_WIDTH `ifdef STREAM42_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM42_OUT_WIDTH , 8'd42 `endif
                `ifdef STREAM43_OUT_WIDTH `ifdef STREAM43_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM43_OUT_WIDTH , 8'd43 `endif
                `ifdef STREAM44_OUT_WIDTH `ifdef STREAM44_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM44_OUT_WIDTH , 8'd44 `endif
                `ifdef STREAM45_OUT_WIDTH `ifdef STREAM45_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM45_OUT_WIDTH , 8'd45 `endif
                `ifdef STREAM46_OUT_WIDTH `ifdef STREAM46_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM46_OUT_WIDTH , 8'd46 `endif
                `ifdef STREAM47_OUT_WIDTH `ifdef STREAM47_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM47_OUT_WIDTH , 8'd47 `endif
                `ifdef STREAM48_OUT_WIDTH `ifdef STREAM48_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM48_OUT_WIDTH , 8'd48 `endif
                `ifdef STREAM49_OUT_WIDTH `ifdef STREAM49_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM49_OUT_WIDTH , 8'd49 `endif
                `ifdef STREAM50_OUT_WIDTH `ifdef STREAM50_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM50_OUT_WIDTH , 8'd50 `endif
                `ifdef STREAM51_OUT_WIDTH `ifdef STREAM51_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM51_OUT_WIDTH , 8'd51 `endif
                `ifdef STREAM52_OUT_WIDTH `ifdef STREAM52_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM52_OUT_WIDTH , 8'd52 `endif
                `ifdef STREAM53_OUT_WIDTH `ifdef STREAM53_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM53_OUT_WIDTH , 8'd53 `endif
                `ifdef STREAM54_OUT_WIDTH `ifdef STREAM54_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM54_OUT_WIDTH , 8'd54 `endif
                `ifdef STREAM55_OUT_WIDTH `ifdef STREAM55_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM55_OUT_WIDTH , 8'd55 `endif
                `ifdef STREAM56_OUT_WIDTH `ifdef STREAM56_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM56_OUT_WIDTH , 8'd56 `endif
                `ifdef STREAM57_OUT_WIDTH `ifdef STREAM57_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM57_OUT_WIDTH , 8'd57 `endif
                `ifdef STREAM58_OUT_WIDTH `ifdef STREAM58_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM58_OUT_WIDTH , 8'd58 `endif
                `ifdef STREAM59_OUT_WIDTH `ifdef STREAM59_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM59_OUT_WIDTH , 8'd59 `endif
                `ifdef STREAM60_OUT_WIDTH `ifdef STREAM60_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM60_OUT_WIDTH , 8'd60 `endif
                `ifdef STREAM61_OUT_WIDTH `ifdef STREAM61_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM61_OUT_WIDTH , 8'd61 `endif
                `ifdef STREAM62_OUT_WIDTH `ifdef STREAM62_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM62_OUT_WIDTH , 8'd62 `endif
                `ifdef STREAM63_OUT_WIDTH `ifdef STREAM63_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM63_OUT_WIDTH , 8'd63 `endif
                `ifdef STREAM64_OUT_WIDTH `ifdef STREAM64_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM64_OUT_WIDTH , 8'd64 `endif
                `ifdef STREAM65_OUT_WIDTH `ifdef STREAM65_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM65_OUT_WIDTH , 8'd65 `endif
                `ifdef STREAM66_OUT_WIDTH `ifdef STREAM66_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM66_OUT_WIDTH , 8'd66 `endif
                `ifdef STREAM67_OUT_WIDTH `ifdef STREAM67_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM67_OUT_WIDTH , 8'd67 `endif
                `ifdef STREAM68_OUT_WIDTH `ifdef STREAM68_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM68_OUT_WIDTH , 8'd68 `endif
                `ifdef STREAM69_OUT_WIDTH `ifdef STREAM69_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM69_OUT_WIDTH , 8'd69 `endif
                `ifdef STREAM70_OUT_WIDTH `ifdef STREAM70_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM70_OUT_WIDTH , 8'd70 `endif
                `ifdef STREAM71_OUT_WIDTH `ifdef STREAM71_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM71_OUT_WIDTH , 8'd71 `endif
                `ifdef STREAM72_OUT_WIDTH `ifdef STREAM72_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM72_OUT_WIDTH , 8'd72 `endif
                `ifdef STREAM73_OUT_WIDTH `ifdef STREAM73_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM73_OUT_WIDTH , 8'd73 `endif
                `ifdef STREAM74_OUT_WIDTH `ifdef STREAM74_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM74_OUT_WIDTH , 8'd74 `endif
                `ifdef STREAM75_OUT_WIDTH `ifdef STREAM75_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM75_OUT_WIDTH , 8'd75 `endif
                `ifdef STREAM76_OUT_WIDTH `ifdef STREAM76_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM76_OUT_WIDTH , 8'd76 `endif
                `ifdef STREAM77_OUT_WIDTH `ifdef STREAM77_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM77_OUT_WIDTH , 8'd77 `endif
                `ifdef STREAM78_OUT_WIDTH `ifdef STREAM78_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM78_OUT_WIDTH , 8'd78 `endif
                `ifdef STREAM79_OUT_WIDTH `ifdef STREAM79_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM79_OUT_WIDTH , 8'd79 `endif
                `ifdef STREAM80_OUT_WIDTH `ifdef STREAM80_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM80_OUT_WIDTH , 8'd80 `endif
                `ifdef STREAM81_OUT_WIDTH `ifdef STREAM81_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM81_OUT_WIDTH , 8'd81 `endif
                `ifdef STREAM82_OUT_WIDTH `ifdef STREAM82_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM82_OUT_WIDTH , 8'd82 `endif
                `ifdef STREAM83_OUT_WIDTH `ifdef STREAM83_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM83_OUT_WIDTH , 8'd83 `endif
                `ifdef STREAM84_OUT_WIDTH `ifdef STREAM84_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM84_OUT_WIDTH , 8'd84 `endif
                `ifdef STREAM85_OUT_WIDTH `ifdef STREAM85_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM85_OUT_WIDTH , 8'd85 `endif
                `ifdef STREAM86_OUT_WIDTH `ifdef STREAM86_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM86_OUT_WIDTH , 8'd86 `endif
                `ifdef STREAM87_OUT_WIDTH `ifdef STREAM87_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM87_OUT_WIDTH , 8'd87 `endif
                `ifdef STREAM88_OUT_WIDTH `ifdef STREAM88_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM88_OUT_WIDTH , 8'd88 `endif
                `ifdef STREAM89_OUT_WIDTH `ifdef STREAM89_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM89_OUT_WIDTH , 8'd89 `endif
                `ifdef STREAM90_OUT_WIDTH `ifdef STREAM90_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM90_OUT_WIDTH , 8'd90 `endif
                `ifdef STREAM91_OUT_WIDTH `ifdef STREAM91_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM91_OUT_WIDTH , 8'd91 `endif
                `ifdef STREAM92_OUT_WIDTH `ifdef STREAM92_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM92_OUT_WIDTH , 8'd92 `endif
                `ifdef STREAM93_OUT_WIDTH `ifdef STREAM93_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM93_OUT_WIDTH , 8'd93 `endif
                `ifdef STREAM94_OUT_WIDTH `ifdef STREAM94_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM94_OUT_WIDTH , 8'd94 `endif
                `ifdef STREAM95_OUT_WIDTH `ifdef STREAM95_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM95_OUT_WIDTH , 8'd95 `endif
                `ifdef STREAM96_OUT_WIDTH `ifdef STREAM96_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM96_OUT_WIDTH , 8'd96 `endif
                `ifdef STREAM97_OUT_WIDTH `ifdef STREAM97_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM97_OUT_WIDTH , 8'd97 `endif
                `ifdef STREAM98_OUT_WIDTH `ifdef STREAM98_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM98_OUT_WIDTH , 8'd98 `endif
                `ifdef STREAM99_OUT_WIDTH `ifdef STREAM99_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM99_OUT_WIDTH , 8'd99 `endif
                `ifdef STREAM100_OUT_WIDTH `ifdef STREAM100_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM100_OUT_WIDTH , 8'd100 `endif
                `ifdef STREAM101_OUT_WIDTH `ifdef STREAM101_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM101_OUT_WIDTH , 8'd101 `endif
                `ifdef STREAM102_OUT_WIDTH `ifdef STREAM102_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM102_OUT_WIDTH , 8'd102 `endif
                `ifdef STREAM103_OUT_WIDTH `ifdef STREAM103_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM103_OUT_WIDTH , 8'd103 `endif
                `ifdef STREAM104_OUT_WIDTH `ifdef STREAM104_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM104_OUT_WIDTH , 8'd104 `endif
                `ifdef STREAM105_OUT_WIDTH `ifdef STREAM105_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM105_OUT_WIDTH , 8'd105 `endif
                `ifdef STREAM106_OUT_WIDTH `ifdef STREAM106_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM106_OUT_WIDTH , 8'd106 `endif
                `ifdef STREAM107_OUT_WIDTH `ifdef STREAM107_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM107_OUT_WIDTH , 8'd107 `endif
                `ifdef STREAM108_OUT_WIDTH `ifdef STREAM108_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM108_OUT_WIDTH , 8'd108 `endif
                `ifdef STREAM109_OUT_WIDTH `ifdef STREAM109_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM109_OUT_WIDTH , 8'd109 `endif
                `ifdef STREAM110_OUT_WIDTH `ifdef STREAM110_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM110_OUT_WIDTH , 8'd110 `endif
                `ifdef STREAM111_OUT_WIDTH `ifdef STREAM111_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM111_OUT_WIDTH , 8'd111 `endif
                `ifdef STREAM112_OUT_WIDTH `ifdef STREAM112_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM112_OUT_WIDTH , 8'd112 `endif
                `ifdef STREAM113_OUT_WIDTH `ifdef STREAM113_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM113_OUT_WIDTH , 8'd113 `endif
                `ifdef STREAM114_OUT_WIDTH `ifdef STREAM114_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM114_OUT_WIDTH , 8'd114 `endif
                `ifdef STREAM115_OUT_WIDTH `ifdef STREAM115_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM115_OUT_WIDTH , 8'd115 `endif
                `ifdef STREAM116_OUT_WIDTH `ifdef STREAM116_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM116_OUT_WIDTH , 8'd116 `endif
                `ifdef STREAM117_OUT_WIDTH `ifdef STREAM117_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM117_OUT_WIDTH , 8'd117 `endif
                `ifdef STREAM118_OUT_WIDTH `ifdef STREAM118_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM118_OUT_WIDTH , 8'd118 `endif
                `ifdef STREAM119_OUT_WIDTH `ifdef STREAM119_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM119_OUT_WIDTH , 8'd119 `endif
                `ifdef STREAM120_OUT_WIDTH `ifdef STREAM120_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM120_OUT_WIDTH , 8'd120 `endif
                `ifdef STREAM121_OUT_WIDTH `ifdef STREAM121_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM121_OUT_WIDTH , 8'd121 `endif
                `ifdef STREAM122_OUT_WIDTH `ifdef STREAM122_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM122_OUT_WIDTH , 8'd122 `endif
                `ifdef STREAM123_OUT_WIDTH `ifdef STREAM123_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM123_OUT_WIDTH , 8'd123 `endif
                `ifdef STREAM124_OUT_WIDTH `ifdef STREAM124_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM124_OUT_WIDTH , 8'd124 `endif
                `ifdef STREAM125_OUT_WIDTH `ifdef STREAM125_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM125_OUT_WIDTH , 8'd125 `endif
                `ifdef STREAM126_OUT_WIDTH `ifdef STREAM126_OUT_256BIT , 32'd2 `else , 32'd1 `endif , 32'd`STREAM126_OUT_WIDTH , 8'd126 `endif
                    };

		`ifndef STREAM1_OUT_256BIT
		   assign stream_out_ow_dvld[1] = 'd1;
		`endif
		`ifndef STREAM2_OUT_256BIT
		   assign stream_out_ow_dvld[2] = 'd1;
		`endif
		`ifndef STREAM3_OUT_256BIT
		   assign stream_out_ow_dvld[3] = 'd1;
		`endif
		`ifndef STREAM4_OUT_256BIT
		   assign stream_out_ow_dvld[4] = 'd1;
		`endif
		`ifndef STREAM5_OUT_256BIT
		   assign stream_out_ow_dvld[5] = 'd1;
		`endif
		`ifndef STREAM6_OUT_256BIT
		   assign stream_out_ow_dvld[6] = 'd1;
		`endif
		`ifndef STREAM7_OUT_256BIT
		   assign stream_out_ow_dvld[7] = 'd1;
		`endif
		`ifndef STREAM8_OUT_256BIT
		   assign stream_out_ow_dvld[8] = 'd1;
		`endif
		`ifndef STREAM9_OUT_256BIT
		   assign stream_out_ow_dvld[9] = 'd1;
		`endif
		`ifndef STREAM10_OUT_256BIT
		   assign stream_out_ow_dvld[10] = 'd1;
		`endif
		`ifndef STREAM11_OUT_256BIT
		   assign stream_out_ow_dvld[11] = 'd1;
		`endif
		`ifndef STREAM12_OUT_256BIT
		   assign stream_out_ow_dvld[12] = 'd1;
		`endif
		`ifndef STREAM13_OUT_256BIT
		   assign stream_out_ow_dvld[13] = 'd1;
		`endif
		`ifndef STREAM14_OUT_256BIT
		   assign stream_out_ow_dvld[14] = 'd1;
		`endif
		`ifndef STREAM15_OUT_256BIT
		   assign stream_out_ow_dvld[15] = 'd1;
		`endif
		`ifndef STREAM16_OUT_256BIT
		   assign stream_out_ow_dvld[16] = 'd1;
		`endif
		`ifndef STREAM17_OUT_256BIT
		   assign stream_out_ow_dvld[17] = 'd1;
		`endif
		`ifndef STREAM18_OUT_256BIT
		   assign stream_out_ow_dvld[18] = 'd1;
		`endif
		`ifndef STREAM19_OUT_256BIT
		   assign stream_out_ow_dvld[19] = 'd1;
		`endif
		`ifndef STREAM20_OUT_256BIT
		   assign stream_out_ow_dvld[20] = 'd1;
		`endif
		`ifndef STREAM21_OUT_256BIT
		   assign stream_out_ow_dvld[21] = 'd1;
		`endif
		`ifndef STREAM22_OUT_256BIT
		   assign stream_out_ow_dvld[22] = 'd1;
		`endif
		`ifndef STREAM23_OUT_256BIT
		   assign stream_out_ow_dvld[23] = 'd1;
		`endif
		`ifndef STREAM24_OUT_256BIT
		   assign stream_out_ow_dvld[24] = 'd1;
		`endif
		`ifndef STREAM25_OUT_256BIT
		   assign stream_out_ow_dvld[25] = 'd1;
		`endif
		`ifndef STREAM26_OUT_256BIT
		   assign stream_out_ow_dvld[26] = 'd1;
		`endif
		`ifndef STREAM27_OUT_256BIT
		   assign stream_out_ow_dvld[27] = 'd1;
		`endif
		`ifndef STREAM28_OUT_256BIT
		   assign stream_out_ow_dvld[28] = 'd1;
		`endif
		`ifndef STREAM29_OUT_256BIT
		   assign stream_out_ow_dvld[29] = 'd1;
		`endif
		`ifndef STREAM30_OUT_256BIT
		   assign stream_out_ow_dvld[30] = 'd1;
		`endif
		`ifndef STREAM31_OUT_256BIT
		   assign stream_out_ow_dvld[31] = 'd1;
		`endif
		`ifndef STREAM32_OUT_256BIT
		   assign stream_out_ow_dvld[32] = 'd1;
		`endif
		`ifndef STREAM33_OUT_256BIT
		   assign stream_out_ow_dvld[33] = 'd1;
		`endif
		`ifndef STREAM34_OUT_256BIT
		   assign stream_out_ow_dvld[34] = 'd1;
		`endif
		`ifndef STREAM35_OUT_256BIT
		   assign stream_out_ow_dvld[35] = 'd1;
		`endif
		`ifndef STREAM36_OUT_256BIT
		   assign stream_out_ow_dvld[36] = 'd1;
		`endif
		`ifndef STREAM37_OUT_256BIT
		   assign stream_out_ow_dvld[37] = 'd1;
		`endif
		`ifndef STREAM38_OUT_256BIT
		   assign stream_out_ow_dvld[38] = 'd1;
		`endif
		`ifndef STREAM39_OUT_256BIT
		   assign stream_out_ow_dvld[39] = 'd1;
		`endif
		`ifndef STREAM40_OUT_256BIT
		   assign stream_out_ow_dvld[40] = 'd1;
		`endif
		`ifndef STREAM41_OUT_256BIT
		   assign stream_out_ow_dvld[41] = 'd1;
		`endif
		`ifndef STREAM42_OUT_256BIT
		   assign stream_out_ow_dvld[42] = 'd1;
		`endif
		`ifndef STREAM43_OUT_256BIT
		   assign stream_out_ow_dvld[43] = 'd1;
		`endif
		`ifndef STREAM44_OUT_256BIT
		   assign stream_out_ow_dvld[44] = 'd1;
		`endif
		`ifndef STREAM45_OUT_256BIT
		   assign stream_out_ow_dvld[45] = 'd1;
		`endif
		`ifndef STREAM46_OUT_256BIT
		   assign stream_out_ow_dvld[46] = 'd1;
		`endif
		`ifndef STREAM47_OUT_256BIT
		   assign stream_out_ow_dvld[47] = 'd1;
		`endif
		`ifndef STREAM48_OUT_256BIT
		   assign stream_out_ow_dvld[48] = 'd1;
		`endif
		`ifndef STREAM49_OUT_256BIT
		   assign stream_out_ow_dvld[49] = 'd1;
		`endif
		`ifndef STREAM50_OUT_256BIT
		   assign stream_out_ow_dvld[50] = 'd1;
		`endif
		`ifndef STREAM51_OUT_256BIT
		   assign stream_out_ow_dvld[51] = 'd1;
		`endif
		`ifndef STREAM52_OUT_256BIT
		   assign stream_out_ow_dvld[52] = 'd1;
		`endif
		`ifndef STREAM53_OUT_256BIT
		   assign stream_out_ow_dvld[53] = 'd1;
		`endif
		`ifndef STREAM54_OUT_256BIT
		   assign stream_out_ow_dvld[54] = 'd1;
		`endif
		`ifndef STREAM55_OUT_256BIT
		   assign stream_out_ow_dvld[55] = 'd1;
		`endif
		`ifndef STREAM56_OUT_256BIT
		   assign stream_out_ow_dvld[56] = 'd1;
		`endif
		`ifndef STREAM57_OUT_256BIT
		   assign stream_out_ow_dvld[57] = 'd1;
		`endif
		`ifndef STREAM58_OUT_256BIT
		   assign stream_out_ow_dvld[58] = 'd1;
		`endif
		`ifndef STREAM59_OUT_256BIT
		   assign stream_out_ow_dvld[59] = 'd1;
		`endif
		`ifndef STREAM60_OUT_256BIT
		   assign stream_out_ow_dvld[60] = 'd1;
		`endif
		`ifndef STREAM61_OUT_256BIT
		   assign stream_out_ow_dvld[61] = 'd1;
		`endif
		`ifndef STREAM62_OUT_256BIT
		   assign stream_out_ow_dvld[62] = 'd1;
		`endif
		`ifndef STREAM63_OUT_256BIT
		   assign stream_out_ow_dvld[63] = 'd1;
		`endif
		`ifndef STREAM64_OUT_256BIT
		   assign stream_out_ow_dvld[64] = 'd1;
		`endif
		`ifndef STREAM65_OUT_256BIT
		   assign stream_out_ow_dvld[65] = 'd1;
		`endif
		`ifndef STREAM66_OUT_256BIT
		   assign stream_out_ow_dvld[66] = 'd1;
		`endif
		`ifndef STREAM67_OUT_256BIT
		   assign stream_out_ow_dvld[67] = 'd1;
		`endif
		`ifndef STREAM68_OUT_256BIT
		   assign stream_out_ow_dvld[68] = 'd1;
		`endif
		`ifndef STREAM69_OUT_256BIT
		   assign stream_out_ow_dvld[69] = 'd1;
		`endif
		`ifndef STREAM70_OUT_256BIT
		   assign stream_out_ow_dvld[70] = 'd1;
		`endif
		`ifndef STREAM71_OUT_256BIT
		   assign stream_out_ow_dvld[71] = 'd1;
		`endif
		`ifndef STREAM72_OUT_256BIT
		   assign stream_out_ow_dvld[72] = 'd1;
		`endif
		`ifndef STREAM73_OUT_256BIT
		   assign stream_out_ow_dvld[73] = 'd1;
		`endif
		`ifndef STREAM74_OUT_256BIT
		   assign stream_out_ow_dvld[74] = 'd1;
		`endif
		`ifndef STREAM75_OUT_256BIT
		   assign stream_out_ow_dvld[75] = 'd1;
		`endif
		`ifndef STREAM76_OUT_256BIT
		   assign stream_out_ow_dvld[76] = 'd1;
		`endif
		`ifndef STREAM77_OUT_256BIT
		   assign stream_out_ow_dvld[77] = 'd1;
		`endif
		`ifndef STREAM78_OUT_256BIT
		   assign stream_out_ow_dvld[78] = 'd1;
		`endif
		`ifndef STREAM79_OUT_256BIT
		   assign stream_out_ow_dvld[79] = 'd1;
		`endif
		`ifndef STREAM80_OUT_256BIT
		   assign stream_out_ow_dvld[80] = 'd1;
		`endif
		`ifndef STREAM81_OUT_256BIT
		   assign stream_out_ow_dvld[81] = 'd1;
		`endif
		`ifndef STREAM82_OUT_256BIT
		   assign stream_out_ow_dvld[82] = 'd1;
		`endif
		`ifndef STREAM83_OUT_256BIT
		   assign stream_out_ow_dvld[83] = 'd1;
		`endif
		`ifndef STREAM84_OUT_256BIT
		   assign stream_out_ow_dvld[84] = 'd1;
		`endif
		`ifndef STREAM85_OUT_256BIT
		   assign stream_out_ow_dvld[85] = 'd1;
		`endif
		`ifndef STREAM86_OUT_256BIT
		   assign stream_out_ow_dvld[86] = 'd1;
		`endif
		`ifndef STREAM87_OUT_256BIT
		   assign stream_out_ow_dvld[87] = 'd1;
		`endif
		`ifndef STREAM88_OUT_256BIT
		   assign stream_out_ow_dvld[88] = 'd1;
		`endif
		`ifndef STREAM89_OUT_256BIT
		   assign stream_out_ow_dvld[89] = 'd1;
		`endif
		`ifndef STREAM90_OUT_256BIT
		   assign stream_out_ow_dvld[90] = 'd1;
		`endif
		`ifndef STREAM91_OUT_256BIT
		   assign stream_out_ow_dvld[91] = 'd1;
		`endif
		`ifndef STREAM92_OUT_256BIT
		   assign stream_out_ow_dvld[92] = 'd1;
		`endif
		`ifndef STREAM93_OUT_256BIT
		   assign stream_out_ow_dvld[93] = 'd1;
		`endif
		`ifndef STREAM94_OUT_256BIT
		   assign stream_out_ow_dvld[94] = 'd1;
		`endif
		`ifndef STREAM95_OUT_256BIT
		   assign stream_out_ow_dvld[95] = 'd1;
		`endif
		`ifndef STREAM96_OUT_256BIT
		   assign stream_out_ow_dvld[96] = 'd1;
		`endif
		`ifndef STREAM97_OUT_256BIT
		   assign stream_out_ow_dvld[97] = 'd1;
		`endif
		`ifndef STREAM98_OUT_256BIT
		   assign stream_out_ow_dvld[98] = 'd1;
		`endif
		`ifndef STREAM99_OUT_256BIT
		   assign stream_out_ow_dvld[99] = 'd1;
		`endif
		`ifndef STREAM100_OUT_256BIT
		   assign stream_out_ow_dvld[100] = 'd1;
		`endif
		`ifndef STREAM101_OUT_256BIT
		   assign stream_out_ow_dvld[101] = 'd1;
		`endif
		`ifndef STREAM102_OUT_256BIT
		   assign stream_out_ow_dvld[102] = 'd1;
		`endif
		`ifndef STREAM103_OUT_256BIT
		   assign stream_out_ow_dvld[103] = 'd1;
		`endif
		`ifndef STREAM104_OUT_256BIT
		   assign stream_out_ow_dvld[104] = 'd1;
		`endif
		`ifndef STREAM105_OUT_256BIT
		   assign stream_out_ow_dvld[105] = 'd1;
		`endif
		`ifndef STREAM106_OUT_256BIT
		   assign stream_out_ow_dvld[106] = 'd1;
		`endif
		`ifndef STREAM107_OUT_256BIT
		   assign stream_out_ow_dvld[107] = 'd1;
		`endif
		`ifndef STREAM108_OUT_256BIT
		   assign stream_out_ow_dvld[108] = 'd1;
		`endif
		`ifndef STREAM109_OUT_256BIT
		   assign stream_out_ow_dvld[109] = 'd1;
		`endif
		`ifndef STREAM110_OUT_256BIT
		   assign stream_out_ow_dvld[110] = 'd1;
		`endif
		`ifndef STREAM111_OUT_256BIT
		   assign stream_out_ow_dvld[111] = 'd1;
		`endif
		`ifndef STREAM112_OUT_256BIT
		   assign stream_out_ow_dvld[112] = 'd1;
		`endif
		`ifndef STREAM113_OUT_256BIT
		   assign stream_out_ow_dvld[113] = 'd1;
		`endif
		`ifndef STREAM114_OUT_256BIT
		   assign stream_out_ow_dvld[114] = 'd1;
		`endif
		`ifndef STREAM115_OUT_256BIT
		   assign stream_out_ow_dvld[115] = 'd1;
		`endif
		`ifndef STREAM116_OUT_256BIT
		   assign stream_out_ow_dvld[116] = 'd1;
		`endif
		`ifndef STREAM117_OUT_256BIT
		   assign stream_out_ow_dvld[117] = 'd1;
		`endif
		`ifndef STREAM118_OUT_256BIT
		   assign stream_out_ow_dvld[118] = 'd1;
		`endif
		`ifndef STREAM119_OUT_256BIT
		   assign stream_out_ow_dvld[119] = 'd1;
		`endif
		`ifndef STREAM120_OUT_256BIT
		   assign stream_out_ow_dvld[120] = 'd1;
		`endif
		`ifndef STREAM121_OUT_256BIT
		   assign stream_out_ow_dvld[121] = 'd1;
		`endif
		`ifndef STREAM122_OUT_256BIT
		   assign stream_out_ow_dvld[122] = 'd1;
		`endif
		`ifndef STREAM123_OUT_256BIT
		   assign stream_out_ow_dvld[123] = 'd1;
		`endif
		`ifndef STREAM124_OUT_256BIT
		   assign stream_out_ow_dvld[124] = 'd1;
		`endif
		`ifndef STREAM125_OUT_256BIT
		   assign stream_out_ow_dvld[125] = 'd1;
		`endif
		`ifndef STREAM126_OUT_256BIT
		   assign stream_out_ow_dvld[126] = 'd1;
		`endif



    genvar k;
    generate
        for( k = 0; |INSTREAM[71+(k*72):0+(k*72)]; k=k+1)
            begin: stream_in
							wire sconv_in_valid, sconv_in_rdy;
							wire [C_DATA_WIDTH-1:0] sconv_in_data;
							wire [OW_DVLD_W-1:0] sconv_in_ow_dvld;
							InStreamWidthConversion #(
									.W(INSTREAM[39+(k*72):8+(k*72)]),
									.C_DATA_WIDTH(C_DATA_WIDTH)
							) gen_width_in (
								.clk(clk),
								.rst(rst),

								.si_valid(sconv_in_valid),
								.si_data(sconv_in_data[C_DATA_WIDTH-1:0]),
								.si_ow_dvld(sconv_in_ow_dvld[OW_DVLD_W-1:0]),
								.si_rdy(sconv_in_rdy),

								.so_valid(stream_in_valid[INSTREAM[7+(k*72):0+(k*72)]]),
								.so_rdy(stream_in_rdy[INSTREAM[7+(k*72):0+(k*72)]]),
								.so_data(stream_in_data[INSTREAM[7+(k*72):0+(k*72)]][INSTREAM[39+(k*72):8+(k*72)]-1:0]),
								.so_ow_dvld(stream_in_ow_dvld[INSTREAM[7+(k*72):0+(k*72)]][INSTREAM[71+(k*72):40+(k*72)]-1:0])
							);
							PicoStreamIn #(
								  .ID(INSTREAM[7+(k*72):0+(k*72)]),
							          .C_DATA_WIDTH(C_DATA_WIDTH)
							 ) gen_stream_in (
								  .clk(clk),
								  .rst(rst),

								  .s_rdy(sconv_in_valid),  //valid
								  .s_en(sconv_in_rdy), // rdy
								  .s_data(sconv_in_data[C_DATA_WIDTH-1:0]),
								  .s_ow_dvld(sconv_in_ow_dvld[OW_DVLD_W-1:0]),

								  .s_in_valid(s_in_valid),
								  .s_in_id(s_in_id[8:0]),
								  .s_in_data(s_in_data[C_DATA_WIDTH-1:0]),
								  .s_in_ow_dvld(s_in_ow_dvld[OW_DVLD_W-1:0]),

								  .s_poll_id(s_poll_id[8:0]),
								  .s_poll_seq(stream_in_desc_poll_seq[INSTREAM[7+(k*72):0+(k*72)]][31:0]),
								  .s_poll_next_desc(stream_in_desc_poll_next_desc[INSTREAM[7+(k*72):0+(k*72)]][127:0]),
								  .s_poll_next_desc_valid(stream_in_desc_poll_next_desc_valid[INSTREAM[7+(k*72):0+(k*72)]]),

								  .s_next_desc_rd_en(s_next_desc_rd_en),
								  .s_next_desc_rd_id(s_next_desc_rd_id[8:0])
							 );
            end
    endgenerate


    `endif //USER_MODULE_NAME


    genvar m;
    generate
        for( m = 0; |OUTSTREAM[71+(m*72):0+(m*72)]; m=m+1)
            begin: stream_out
							wire sconv_out_valid, sconv_out_rdy;
							wire [C_DATA_WIDTH-1:0] sconv_out_data;
							wire [OW_DVLD_W-1:0] sconv_out_ow_dvld;
							OutStreamWidthConversion #(
									.W(OUTSTREAM[39+(m*72):8+(m*72)]),
									.C_DATA_WIDTH(C_DATA_WIDTH)
							) gen_width_out (
								.clk(clk),
								.rst(rst),

								.so_valid(sconv_out_valid),
								.so_data(sconv_out_data[C_DATA_WIDTH-1:0]),
								.so_ow_dvld(sconv_out_ow_dvld[OW_DVLD_W-1:0]),
								.so_rdy(sconv_out_rdy),

								.si_valid(stream_out_valid[OUTSTREAM[7+(m*72):0+(m*72)]]),
								.si_rdy(stream_out_rdy[OUTSTREAM[7+(m*72):0+(m*72)]]),
								.si_data(stream_out_data[OUTSTREAM[7+(m*72):0+(m*72)]][OUTSTREAM[39+(m*72):8+(m*72)]-1:0]),
								.si_ow_dvld(stream_out_ow_dvld[OUTSTREAM[7+(m*72):0+(m*72)]][OUTSTREAM[71+(m*72):40+(m*72)]-1:0])
							);

							PicoStreamOut #(
							  .ID(OUTSTREAM[7+(m*72):0+(m*72)]),
							  .C_DATA_WIDTH(C_DATA_WIDTH)
							) gen_stream_out (
							  .clk(clk),
							  .rst(rst),

							  .s_rdy(sconv_out_rdy),
							  .s_valid(sconv_out_valid),
							  .s_data(sconv_out_data[C_DATA_WIDTH-1:0]),
							  .s_ow_dvld(sconv_out_ow_dvld[OW_DVLD_W-1:0]),

							  .s_out_en(s_out_en),
							  .s_out_id(s_out_id[8:0]),
							  .s_out_data(stream_out_data_card[OUTSTREAM[7+(m*72):0+(m*72)]][C_DATA_WIDTH-1:0]),
							  .s_out_ow_dvld(stream_out_ow_dvld_card[OUTSTREAM[7+(m*72):0+(m*72)]][OW_DVLD_W-1:0]),

							  .s_in_valid(s_in_valid),
							  .s_in_id(s_in_id[8:0]),
							  .s_in_data(s_in_data[C_DATA_WIDTH-1:0]),
							  .s_in_ow_dvld(s_in_ow_dvld[OW_DVLD_W-1:0]),

							  .s_poll_id(s_poll_id[8:0]),
							  .s_poll_seq(stream_out_desc_poll_seq[OUTSTREAM[7+(m*72):0+(m*72)]][31:0]),
							  .s_poll_next_desc(stream_out_desc_poll_next_desc[OUTSTREAM[7+(m*72):0+(m*72)]][127:0]),
							  .s_poll_next_desc_valid(stream_out_desc_poll_next_desc_valid[OUTSTREAM[7+(m*72):0+(m*72)]]),

							  .s_next_desc_rd_en(s_next_desc_rd_en),
							  .s_next_desc_rd_id(s_next_desc_rd_id[8:0])
						 );
            end
    endgenerate

    // end usermodule stream interface

`ifdef USER_MODULE_NAME
    `USER_MODULE_NAME
      `ifdef PICO_DDR3_OR_DDR4
         #(
            .C0_C_S_AXI_ID_WIDTH       ( C0_C_S_AXI_ID_WIDTH-4 ),
            .C0_C_S_AXI_ADDR_WIDTH     ( C0_C_S_AXI_ADDR_WIDTH ),
            .C0_C_S_AXI_DATA_WIDTH     ( C0_C_S_AXI_DATA_WIDTH )
         )
      `endif // PICO_DDR3_OR_DDR4
     UserModule (
    `undef UM_PREPEND_COMMA      // In case this gets used before
    `undef INCLUDE_STREAM_COMMON // ditto

    `ifdef EXTRA_CLK
         `ifdef  UM_PREPEND_COMMA , `endif
         `define UM_PREPEND_COMMA
         .extra_clk(extra_clk)
    `endif

    `ifdef USER_DIRECT_PCI
         `ifdef  UM_PREPEND_COMMA , `endif
         `define UM_PREPEND_COMMA
        .user_pci_wr_q_data(user_pci_wr_q_data),
        .user_pci_wr_q_valid(user_pci_wr_q_valid),
        .user_pci_wr_q_en(user_pci_wr_q_en),

        .user_pci_wr_data_q_data(user_pci_wr_data_q_data),
        .user_pci_wr_data_q_valid(user_pci_wr_data_q_valid),
        .user_pci_wr_data_q_en(user_pci_wr_data_q_en),

        .direct_rx_valid(direct_rx_valid),
        .direct_rx_data(s_in_data[C_DATA_WIDTH-1:0])
    `endif

    `ifdef PICOBUS_WIDTH
         `ifdef  UM_PREPEND_COMMA , `endif
         `define UM_PREPEND_COMMA
        .PicoClk(UserModulePicoClk),
        .PicoRst(UserModulePicoRst),
        .PicoAddr(UserModulePicoAddr[31:0]),
        .PicoDataIn(UserModulePicoDataIn),
        .PicoRd(UserModulePicoRd),
        .PicoWr(UserModulePicoWr),
        .PicoDataOut(UserModulePicoDataOut)
    `endif

`ifdef ENABLE_HMC
         `ifdef  UM_PREPEND_COMMA , `endif
         `define UM_PREPEND_COMMA
    `ifdef USE_512_BIT_HMC_CONTROLLER
        .hmc_clk_p0                   ( hmc_axi_port[0].clk     ) ,


        .axi_awid_p0                  ( hmc_axi_port[0].awid    ) ,
        .axi_awaddr_p0                ( hmc_axi_port[0].awaddr  ) ,
        .axi_awlen_p0                 ( hmc_axi_port[0].awlen   ) ,
        .axi_awsize_p0                ( hmc_axi_port[0].awsize  ) ,
        .axi_awburst_p0               ( hmc_axi_port[0].awburst ) ,
        .axi_awlock_p0                ( hmc_axi_port[0].awlock  ) ,
        .axi_awcache_p0               ( hmc_axi_port[0].awcache ) ,
        .axi_awprot_p0                ( hmc_axi_port[0].awprot  ) ,
        .axi_awqos_p0                 ( hmc_axi_port[0].awqos   ) ,
        .axi_awvalid_p0               ( hmc_axi_port[0].awvalid ) ,
        .axi_awready_p0               ( hmc_axi_port[0].awready ) ,
        .axi_wdata_p0                 ( hmc_axi_port[0].wdata   ) ,

        .axi_wstrb_p0                 ( hmc_axi_port[0].wstrb   ) ,
        .axi_wlast_p0                 ( hmc_axi_port[0].wlast   ) ,
        .axi_wvalid_p0                ( hmc_axi_port[0].wvalid  ) ,
        .axi_wready_p0                ( hmc_axi_port[0].wready  ) ,
        .axi_bid_p0                   ( hmc_axi_port[0].bid     ) ,
        .axi_bresp_p0                 ( hmc_axi_port[0].bresp   ) ,
        .axi_bvalid_p0                ( hmc_axi_port[0].bvalid  ) ,
        .axi_bready_p0                ( hmc_axi_port[0].bready  ) ,
        .axi_arid_p0                  ( hmc_axi_port[0].arid    ) ,
        .axi_araddr_p0                ( hmc_axi_port[0].araddr  ) ,
        .axi_arlen_p0                 ( hmc_axi_port[0].arlen   ) ,
        .axi_arsize_p0                ( hmc_axi_port[0].arsize  ) ,
        .axi_arburst_p0               ( hmc_axi_port[0].arburst ) ,
        .axi_arlock_p0                ( hmc_axi_port[0].arlock  ) ,
        .axi_arcache_p0               ( hmc_axi_port[0].arcache ) ,
        .axi_arprot_p0                ( hmc_axi_port[0].arprot  ) ,
        .axi_arqos_p0                 ( hmc_axi_port[0].arqos   ) ,
        .axi_arvalid_p0               ( hmc_axi_port[0].arvalid ) ,
        .axi_arready_p0               ( hmc_axi_port[0].arready ) ,
        .axi_rid_p0                   ( hmc_axi_port[0].rid     ) ,
        .axi_rdata_p0                 ( hmc_axi_port[0].rdata   ) ,
        .axi_rresp_p0                 ( hmc_axi_port[0].rresp   ) ,
        .axi_rlast_p0                 ( hmc_axi_port[0].rlast   ) ,
        .axi_rvalid_p0                ( hmc_axi_port[0].rvalid  ) ,
        .axi_rready_p0                ( hmc_axi_port[0].rready  ) ,

        .axi_wid_p0                   ( hmc_axi_port[0].wid        ),
        .axi_stride_num_p0            ( hmc_axi_port[0].stride_num ),
        .axi_stride_p0                ( hmc_axi_port[0].stride     ),
        .tags_almostempty_p0          ( hmc_axi_port[0].tags_almostempty ) ,

      `ifdef ENABLE_2ND_HMC_LINK
        // 128-bit port, second controller
        .hmc_clk_p1                      ( hmc_port[1].clk ),
        .hmc_addr_p1                     ( hmc_port[1].addr ),
        .hmc_size_p1                     ( hmc_port[1].size ),
        .hmc_tag_p1                      ( hmc_port[1].tag ),
        .hmc_cmd_valid_p1                ( hmc_port[1].cmd_valid ),
        .hmc_cmd_ready_p1                ( hmc_port[1].cmd_ready ),
        .hmc_cmd_p1                      ( hmc_port[1].cmd ),
        .hmc_wr_data_p1                  ( hmc_port[1].wr_data ),
        .hmc_wr_data_valid_p1            ( hmc_port[1].wr_data_valid ),
        .hmc_wr_data_ready_p1            ( hmc_port[1].wr_data_ready ),
        .hmc_rd_data_p1                  ( hmc_port[1].rd_data ),
        .hmc_rd_data_tag_p1              ( hmc_port[1].rd_data_tag ),
        .hmc_rd_data_valid_p1            ( hmc_port[1].rd_data_valid ),
        .hmc_errstat_p1                  ( hmc_port[1].errstat ),
        .hmc_dinv_p1                     ( hmc_port[1].dinv ),

        // 512-bit AXI port, second controller
        .hmc_clk_p2                   ( hmc_axi_port[1].clk     ) ,


        .axi_awid_p2                  ( hmc_axi_port[1].awid    ) ,
        .axi_awaddr_p2                ( hmc_axi_port[1].awaddr  ) ,
        .axi_awlen_p2                 ( hmc_axi_port[1].awlen   ) ,
        .axi_awsize_p2                ( hmc_axi_port[1].awsize  ) ,
        .axi_awburst_p2               ( hmc_axi_port[1].awburst ) ,
        .axi_awlock_p2                ( hmc_axi_port[1].awlock  ) ,
        .axi_awcache_p2               ( hmc_axi_port[1].awcache ) ,
        .axi_awprot_p2                ( hmc_axi_port[1].awprot  ) ,
        .axi_awqos_p2                 ( hmc_axi_port[1].awqos   ) ,
        .axi_awvalid_p2               ( hmc_axi_port[1].awvalid ) ,
        .axi_awready_p2               ( hmc_axi_port[1].awready ) ,
        .axi_wdata_p2                 ( hmc_axi_port[1].wdata   ) ,

        .axi_wstrb_p2                 ( hmc_axi_port[1].wstrb   ) ,
        .axi_wlast_p2                 ( hmc_axi_port[1].wlast   ) ,
        .axi_wvalid_p2                ( hmc_axi_port[1].wvalid  ) ,
        .axi_wready_p2                ( hmc_axi_port[1].wready  ) ,
        .axi_bid_p2                   ( hmc_axi_port[1].bid     ) ,
        .axi_bresp_p2                 ( hmc_axi_port[1].bresp   ) ,
        .axi_bvalid_p2                ( hmc_axi_port[1].bvalid  ) ,
        .axi_bready_p2                ( hmc_axi_port[1].bready  ) ,
        .axi_arid_p2                  ( hmc_axi_port[1].arid    ) ,
        .axi_araddr_p2                ( hmc_axi_port[1].araddr  ) ,
        .axi_arlen_p2                 ( hmc_axi_port[1].arlen   ) ,
        .axi_arsize_p2                ( hmc_axi_port[1].arsize  ) ,
        .axi_arburst_p2               ( hmc_axi_port[1].arburst ) ,
        .axi_arlock_p2                ( hmc_axi_port[1].arlock  ) ,
        .axi_arcache_p2               ( hmc_axi_port[1].arcache ) ,
        .axi_arprot_p2                ( hmc_axi_port[1].arprot  ) ,
        .axi_arqos_p2                 ( hmc_axi_port[1].arqos   ) ,
        .axi_arvalid_p2               ( hmc_axi_port[1].arvalid ) ,
        .axi_arready_p2               ( hmc_axi_port[1].arready ) ,
        .axi_rid_p2                   ( hmc_axi_port[1].rid     ) ,
        .axi_rdata_p2                 ( hmc_axi_port[1].rdata   ) ,
        .axi_rresp_p2                 ( hmc_axi_port[1].rresp   ) ,
        .axi_rlast_p2                 ( hmc_axi_port[1].rlast   ) ,
        .axi_rvalid_p2                ( hmc_axi_port[1].rvalid  ) ,
        .axi_rready_p2                ( hmc_axi_port[1].rready  ) ,

        .axi_wid_p2                   ( hmc_axi_port[1].wid        ),
        .axi_stride_num_p2            ( hmc_axi_port[1].stride_num ),
        .axi_stride_p2                ( hmc_axi_port[1].stride     ),
        .tags_almostempty_p2          ( hmc_axi_port[1].tags_almostempty ) ,
      `endif // ENABLE_2ND_HMC_LINK

      `ifdef ENABLE_3RD_HMC_LINK
        .hmc_clk_p3                      ( hmc_port[2].clk ),
        .hmc_addr_p3                     ( hmc_port[2].addr ),
        .hmc_size_p3                     ( hmc_port[2].size ),
        .hmc_tag_p3                      ( hmc_port[2].tag ),
        .hmc_cmd_valid_p3                ( hmc_port[2].cmd_valid ),
        .hmc_cmd_ready_p3                ( hmc_port[2].cmd_ready ),
        .hmc_cmd_p3                      ( hmc_port[2].cmd ),
        .hmc_wr_data_p3                  ( hmc_port[2].wr_data ),
        .hmc_wr_data_valid_p3            ( hmc_port[2].wr_data_valid ),
        .hmc_wr_data_ready_p3            ( hmc_port[2].wr_data_ready ),
        .hmc_rd_data_p3                  ( hmc_port[2].rd_data ),
        .hmc_rd_data_tag_p3              ( hmc_port[2].rd_data_tag ),
        .hmc_rd_data_valid_p3            ( hmc_port[2].rd_data_valid ),
        .hmc_errstat_p3                  ( hmc_port[2].errstat ),
        .hmc_dinv_p3                     ( hmc_port[2].dinv ),

        // 512-bit AXI port
        .hmc_clk_p4                   ( hmc_axi_port[2].clk     ) ,


        .axi_awid_p4                  ( hmc_axi_port[2].awid    ) ,
        .axi_awaddr_p4                ( hmc_axi_port[2].awaddr  ) ,
        .axi_awlen_p4                 ( hmc_axi_port[2].awlen   ) ,
        .axi_awsize_p4                ( hmc_axi_port[2].awsize  ) ,
        .axi_awburst_p4               ( hmc_axi_port[2].awburst ) ,
        .axi_awlock_p4                ( hmc_axi_port[2].awlock  ) ,
        .axi_awcache_p4               ( hmc_axi_port[2].awcache ) ,
        .axi_awprot_p4                ( hmc_axi_port[2].awprot  ) ,
        .axi_awqos_p4                 ( hmc_axi_port[2].awqos   ) ,
        .axi_awvalid_p4               ( hmc_axi_port[2].awvalid ) ,
        .axi_awready_p4               ( hmc_axi_port[2].awready ) ,
        .axi_wdata_p4                 ( hmc_axi_port[2].wdata   ) ,

        .axi_wstrb_p4                 ( hmc_axi_port[2].wstrb   ) ,
        .axi_wlast_p4                 ( hmc_axi_port[2].wlast   ) ,
        .axi_wvalid_p4                ( hmc_axi_port[2].wvalid  ) ,
        .axi_wready_p4                ( hmc_axi_port[2].wready  ) ,
        .axi_bid_p4                   ( hmc_axi_port[2].bid     ) ,
        .axi_bresp_p4                 ( hmc_axi_port[2].bresp   ) ,
        .axi_bvalid_p4                ( hmc_axi_port[2].bvalid  ) ,
        .axi_bready_p4                ( hmc_axi_port[2].bready  ) ,
        .axi_arid_p4                  ( hmc_axi_port[2].arid    ) ,
        .axi_araddr_p4                ( hmc_axi_port[2].araddr  ) ,
        .axi_arlen_p4                 ( hmc_axi_port[2].arlen   ) ,
        .axi_arsize_p4                ( hmc_axi_port[2].arsize  ) ,
        .axi_arburst_p4               ( hmc_axi_port[2].arburst ) ,
        .axi_arlock_p4                ( hmc_axi_port[2].arlock  ) ,
        .axi_arcache_p4               ( hmc_axi_port[2].arcache ) ,
        .axi_arprot_p4                ( hmc_axi_port[2].arprot  ) ,
        .axi_arqos_p4                 ( hmc_axi_port[2].arqos   ) ,
        .axi_arvalid_p4               ( hmc_axi_port[2].arvalid ) ,
        .axi_arready_p4               ( hmc_axi_port[2].arready ) ,
        .axi_rid_p4                   ( hmc_axi_port[2].rid     ) ,
        .axi_rdata_p4                 ( hmc_axi_port[2].rdata   ) ,
        .axi_rresp_p4                 ( hmc_axi_port[2].rresp   ) ,
        .axi_rlast_p4                 ( hmc_axi_port[2].rlast   ) ,
        .axi_rvalid_p4                ( hmc_axi_port[2].rvalid  ) ,
        .axi_rready_p4                ( hmc_axi_port[2].rready  ) ,

        .axi_wid_p4                   ( hmc_axi_port[2].wid        ),
        .axi_stride_num_p4            ( hmc_axi_port[2].stride_num ),
        .axi_stride_p4                ( hmc_axi_port[2].stride     ),
        .tags_almostempty_p4          ( hmc_axi_port[2].tags_almostempty ) ,
      `endif // ENABLE_3RD_HMC_LINK


      `ifdef ENABLE_4TH_HMC_LINK
        .hmc_clk_p5                      ( hmc_port[3].clk ),
        .hmc_addr_p5                     ( hmc_port[3].addr ),
        .hmc_size_p5                     ( hmc_port[3].size ),
        .hmc_tag_p5                      ( hmc_port[3].tag ),
        .hmc_cmd_valid_p5                ( hmc_port[3].cmd_valid ),
        .hmc_cmd_ready_p5                ( hmc_port[3].cmd_ready ),
        .hmc_cmd_p5                      ( hmc_port[3].cmd ),
        .hmc_wr_data_p5                  ( hmc_port[3].wr_data ),
        .hmc_wr_data_valid_p5            ( hmc_port[3].wr_data_valid ),
        .hmc_wr_data_ready_p5            ( hmc_port[3].wr_data_ready ),
        .hmc_rd_data_p5                  ( hmc_port[3].rd_data ),
        .hmc_rd_data_tag_p5              ( hmc_port[3].rd_data_tag ),
        .hmc_rd_data_valid_p5            ( hmc_port[3].rd_data_valid ),
        .hmc_errstat_p5                  ( hmc_port[3].errstat ),
        .hmc_dinv_p5                     ( hmc_port[3].dinv ),

        // 512-bit AXI port
        .hmc_clk_p6                   ( hmc_axi_port[3].clk     ) ,


        .axi_awid_p6                  ( hmc_axi_port[3].awid    ) ,
        .axi_awaddr_p6                ( hmc_axi_port[3].awaddr  ) ,
        .axi_awlen_p6                 ( hmc_axi_port[3].awlen   ) ,
        .axi_awsize_p6                ( hmc_axi_port[3].awsize  ) ,
        .axi_awburst_p6               ( hmc_axi_port[3].awburst ) ,
        .axi_awlock_p6                ( hmc_axi_port[3].awlock  ) ,
        .axi_awcache_p6               ( hmc_axi_port[3].awcache ) ,
        .axi_awprot_p6                ( hmc_axi_port[3].awprot  ) ,
        .axi_awqos_p6                 ( hmc_axi_port[3].awqos   ) ,
        .axi_awvalid_p6               ( hmc_axi_port[3].awvalid ) ,
        .axi_awready_p6               ( hmc_axi_port[3].awready ) ,
        .axi_wdata_p6                 ( hmc_axi_port[3].wdata   ) ,

        .axi_wstrb_p6                 ( hmc_axi_port[3].wstrb   ) ,
        .axi_wlast_p6                 ( hmc_axi_port[3].wlast   ) ,
        .axi_wvalid_p6                ( hmc_axi_port[3].wvalid  ) ,
        .axi_wready_p6                ( hmc_axi_port[3].wready  ) ,
        .axi_bid_p6                   ( hmc_axi_port[3].bid     ) ,
        .axi_bresp_p6                 ( hmc_axi_port[3].bresp   ) ,
        .axi_bvalid_p6                ( hmc_axi_port[3].bvalid  ) ,
        .axi_bready_p6                ( hmc_axi_port[3].bready  ) ,
        .axi_arid_p6                  ( hmc_axi_port[3].arid    ) ,
        .axi_araddr_p6                ( hmc_axi_port[3].araddr  ) ,
        .axi_arlen_p6                 ( hmc_axi_port[3].arlen   ) ,
        .axi_arsize_p6                ( hmc_axi_port[3].arsize  ) ,
        .axi_arburst_p6               ( hmc_axi_port[3].arburst ) ,
        .axi_arlock_p6                ( hmc_axi_port[3].arlock  ) ,
        .axi_arcache_p6               ( hmc_axi_port[3].arcache ) ,
        .axi_arprot_p6                ( hmc_axi_port[3].arprot  ) ,
        .axi_arqos_p6                 ( hmc_axi_port[3].arqos   ) ,
        .axi_arvalid_p6               ( hmc_axi_port[3].arvalid ) ,
        .axi_arready_p6               ( hmc_axi_port[3].arready ) ,
        .axi_rid_p6                   ( hmc_axi_port[3].rid     ) ,
        .axi_rdata_p6                 ( hmc_axi_port[3].rdata   ) ,
        .axi_rresp_p6                 ( hmc_axi_port[3].rresp   ) ,
        .axi_rlast_p6                 ( hmc_axi_port[3].rlast   ) ,
        .axi_rvalid_p6                ( hmc_axi_port[3].rvalid  ) ,
        .axi_rready_p6                ( hmc_axi_port[3].rready  ) ,

        .axi_wid_p6                   ( hmc_axi_port[3].wid        ),
        .axi_stride_num_p6            ( hmc_axi_port[3].stride_num ),
        .axi_stride_p6                ( hmc_axi_port[3].stride     ),
        .tags_almostempty_p6          ( hmc_axi_port[3].tags_almostempty ) ,
      `endif // ENABLE_4TH_HMC_LINK

    `else //USE_512_BIT_HMC_CONTROLLER
        .hmc_clk_p0                      ( hmc_port[1].clk ),
        .hmc_addr_p0                     ( hmc_port[1].addr ),
        .hmc_size_p0                     ( hmc_port[1].size ),
        .hmc_tag_p0                      ( hmc_port[1].tag ),
        .hmc_cmd_valid_p0                ( hmc_port[1].cmd_valid ),
        .hmc_cmd_ready_p0                ( hmc_port[1].cmd_ready ),
        .hmc_cmd_p0                      ( hmc_port[1].cmd ),
        .hmc_wr_data_p0                  ( hmc_port[1].wr_data ),
        .hmc_wr_data_valid_p0            ( hmc_port[1].wr_data_valid ),
        .hmc_wr_data_ready_p0            ( hmc_port[1].wr_data_ready ),
        .hmc_rd_data_p0                  ( hmc_port[1].rd_data ),
        .hmc_rd_data_tag_p0              ( hmc_port[1].rd_data_tag ),
        .hmc_rd_data_valid_p0            ( hmc_port[1].rd_data_valid ),
        .hmc_errstat_p0                  ( hmc_port[1].errstat ),
        .hmc_dinv_p0                     ( hmc_port[1].dinv ),
        .hmc_clk_p1                      ( hmc_port[2].clk ),
        .hmc_addr_p1                     ( hmc_port[2].addr ),
        .hmc_size_p1                     ( hmc_port[2].size ),
        .hmc_tag_p1                      ( hmc_port[2].tag ),
        .hmc_cmd_valid_p1                ( hmc_port[2].cmd_valid ),
        .hmc_cmd_ready_p1                ( hmc_port[2].cmd_ready ),
        .hmc_cmd_p1                      ( hmc_port[2].cmd ),
        .hmc_wr_data_p1                  ( hmc_port[2].wr_data ),
        .hmc_wr_data_valid_p1            ( hmc_port[2].wr_data_valid ),
        .hmc_wr_data_ready_p1            ( hmc_port[2].wr_data_ready ),
        .hmc_rd_data_p1                  ( hmc_port[2].rd_data ),
        .hmc_rd_data_tag_p1              ( hmc_port[2].rd_data_tag ),
        .hmc_rd_data_valid_p1            ( hmc_port[2].rd_data_valid ),
        .hmc_errstat_p1                  ( hmc_port[2].errstat ),
        .hmc_dinv_p1                     ( hmc_port[2].dinv ),
        .hmc_clk_p2                      ( hmc_port[3].clk ),
        .hmc_addr_p2                     ( hmc_port[3].addr ),
        .hmc_size_p2                     ( hmc_port[3].size ),
        .hmc_tag_p2                      ( hmc_port[3].tag ),
        .hmc_cmd_valid_p2                ( hmc_port[3].cmd_valid ),
        .hmc_cmd_ready_p2                ( hmc_port[3].cmd_ready ),
        .hmc_cmd_p2                      ( hmc_port[3].cmd ),
        .hmc_wr_data_p2                  ( hmc_port[3].wr_data ),
        .hmc_wr_data_valid_p2            ( hmc_port[3].wr_data_valid ),
        .hmc_wr_data_ready_p2            ( hmc_port[3].wr_data_ready ),
        .hmc_rd_data_p2                  ( hmc_port[3].rd_data ),
        .hmc_rd_data_tag_p2              ( hmc_port[3].rd_data_tag ),
        .hmc_rd_data_valid_p2            ( hmc_port[3].rd_data_valid ),
        .hmc_errstat_p2                  ( hmc_port[3].errstat ),
        .hmc_dinv_p2                     ( hmc_port[3].dinv ),
        .hmc_clk_p3                      ( hmc_port[4].clk ),
        .hmc_addr_p3                     ( hmc_port[4].addr ),
        .hmc_size_p3                     ( hmc_port[4].size ),
        .hmc_tag_p3                      ( hmc_port[4].tag ),
        .hmc_cmd_valid_p3                ( hmc_port[4].cmd_valid ),
        .hmc_cmd_ready_p3                ( hmc_port[4].cmd_ready ),
        .hmc_cmd_p3                      ( hmc_port[4].cmd ),
        .hmc_wr_data_p3                  ( hmc_port[4].wr_data ),
        .hmc_wr_data_valid_p3            ( hmc_port[4].wr_data_valid ),
        .hmc_wr_data_ready_p3            ( hmc_port[4].wr_data_ready ),
        .hmc_rd_data_p3                  ( hmc_port[4].rd_data ),
        .hmc_rd_data_tag_p3              ( hmc_port[4].rd_data_tag ),
        .hmc_rd_data_valid_p3            ( hmc_port[4].rd_data_valid ),
        .hmc_errstat_p3                  ( hmc_port[4].errstat ),
        .hmc_dinv_p3                     ( hmc_port[4].dinv ),
      `ifdef ENABLE_2ND_HMC_LINK
        .hmc_clk_p4                      ( hmc_port[5].clk ),
        .hmc_addr_p4                     ( hmc_port[5].addr ),
        .hmc_size_p4                     ( hmc_port[5].size ),
        .hmc_tag_p4                      ( hmc_port[5].tag ),
        .hmc_cmd_valid_p4                ( hmc_port[5].cmd_valid ),
        .hmc_cmd_ready_p4                ( hmc_port[5].cmd_ready ),
        .hmc_cmd_p4                      ( hmc_port[5].cmd ),
        .hmc_wr_data_p4                  ( hmc_port[5].wr_data ),
        .hmc_wr_data_valid_p4            ( hmc_port[5].wr_data_valid ),
        .hmc_wr_data_ready_p4            ( hmc_port[5].wr_data_ready ),
        .hmc_rd_data_p4                  ( hmc_port[5].rd_data ),
        .hmc_rd_data_tag_p4              ( hmc_port[5].rd_data_tag ),
        .hmc_rd_data_valid_p4            ( hmc_port[5].rd_data_valid ),
        .hmc_errstat_p4                  ( hmc_port[5].errstat ),
        .hmc_dinv_p4                     ( hmc_port[5].dinv ),
        .hmc_clk_p5                      ( hmc_port[6].clk ),
        .hmc_addr_p5                     ( hmc_port[6].addr ),
        .hmc_size_p5                     ( hmc_port[6].size ),
        .hmc_tag_p5                      ( hmc_port[6].tag ),
        .hmc_cmd_valid_p5                ( hmc_port[6].cmd_valid ),
        .hmc_cmd_ready_p5                ( hmc_port[6].cmd_ready ),
        .hmc_cmd_p5                      ( hmc_port[6].cmd ),
        .hmc_wr_data_p5                  ( hmc_port[6].wr_data ),
        .hmc_wr_data_valid_p5            ( hmc_port[6].wr_data_valid ),
        .hmc_wr_data_ready_p5            ( hmc_port[6].wr_data_ready ),
        .hmc_rd_data_p5                  ( hmc_port[6].rd_data ),
        .hmc_rd_data_tag_p5              ( hmc_port[6].rd_data_tag ),
        .hmc_rd_data_valid_p5            ( hmc_port[6].rd_data_valid ),
        .hmc_errstat_p5                  ( hmc_port[6].errstat ),
        .hmc_dinv_p5                     ( hmc_port[6].dinv ),
        .hmc_clk_p6                      ( hmc_port[7].clk ),
        .hmc_addr_p6                     ( hmc_port[7].addr ),
        .hmc_size_p6                     ( hmc_port[7].size ),
        .hmc_tag_p6                      ( hmc_port[7].tag ),
        .hmc_cmd_valid_p6                ( hmc_port[7].cmd_valid ),
        .hmc_cmd_ready_p6                ( hmc_port[7].cmd_ready ),
        .hmc_cmd_p6                      ( hmc_port[7].cmd ),
        .hmc_wr_data_p6                  ( hmc_port[7].wr_data ),
        .hmc_wr_data_valid_p6            ( hmc_port[7].wr_data_valid ),
        .hmc_wr_data_ready_p6            ( hmc_port[7].wr_data_ready ),
        .hmc_rd_data_p6                  ( hmc_port[7].rd_data ),
        .hmc_rd_data_tag_p6              ( hmc_port[7].rd_data_tag ),
        .hmc_rd_data_valid_p6            ( hmc_port[7].rd_data_valid ),
        .hmc_errstat_p6                  ( hmc_port[7].errstat ),
        .hmc_dinv_p6                     ( hmc_port[7].dinv ),
        .hmc_clk_p7                      ( hmc_port[8].clk ),
        .hmc_addr_p7                     ( hmc_port[8].addr ),
        .hmc_size_p7                     ( hmc_port[8].size ),
        .hmc_tag_p7                      ( hmc_port[8].tag ),
        .hmc_cmd_valid_p7                ( hmc_port[8].cmd_valid ),
        .hmc_cmd_ready_p7                ( hmc_port[8].cmd_ready ),
        .hmc_cmd_p7                      ( hmc_port[8].cmd ),
        .hmc_wr_data_p7                  ( hmc_port[8].wr_data ),
        .hmc_wr_data_valid_p7            ( hmc_port[8].wr_data_valid ),
        .hmc_wr_data_ready_p7            ( hmc_port[8].wr_data_ready ),
        .hmc_rd_data_p7                  ( hmc_port[8].rd_data ),
        .hmc_rd_data_tag_p7              ( hmc_port[8].rd_data_tag ),
        .hmc_rd_data_valid_p7            ( hmc_port[8].rd_data_valid ),
        .hmc_errstat_p7                  ( hmc_port[8].errstat ),
        .hmc_dinv_p7                     ( hmc_port[8].dinv ),
        .hmc_clk_p8                      ( hmc_port[9].clk ),
        .hmc_addr_p8                     ( hmc_port[9].addr ),
        .hmc_size_p8                     ( hmc_port[9].size ),
        .hmc_tag_p8                      ( hmc_port[9].tag ),
        .hmc_cmd_valid_p8                ( hmc_port[9].cmd_valid ),
        .hmc_cmd_ready_p8                ( hmc_port[9].cmd_ready ),
        .hmc_cmd_p8                      ( hmc_port[9].cmd ),
        .hmc_wr_data_p8                  ( hmc_port[9].wr_data ),
        .hmc_wr_data_valid_p8            ( hmc_port[9].wr_data_valid ),
        .hmc_wr_data_ready_p8            ( hmc_port[9].wr_data_ready ),
        .hmc_rd_data_p8                  ( hmc_port[9].rd_data ),
        .hmc_rd_data_tag_p8              ( hmc_port[9].rd_data_tag ),
        .hmc_rd_data_valid_p8            ( hmc_port[9].rd_data_valid ),
        .hmc_errstat_p8                  ( hmc_port[9].errstat ),
        .hmc_dinv_p8                     ( hmc_port[9].dinv ),
	  `endif // ENABLE_2ND_HMC_LINK
      `ifdef ENABLE_3RD_HMC_LINK
        .hmc_clk_p9                      ( hmc_port[10].clk ),
        .hmc_addr_p9                     ( hmc_port[10].addr ),
        .hmc_size_p9                     ( hmc_port[10].size ),
        .hmc_tag_p9                      ( hmc_port[10].tag ),
        .hmc_cmd_valid_p9                ( hmc_port[10].cmd_valid ),
        .hmc_cmd_ready_p9                ( hmc_port[10].cmd_ready ),
        .hmc_cmd_p9                      ( hmc_port[10].cmd ),
        .hmc_wr_data_p9                  ( hmc_port[10].wr_data ),
        .hmc_wr_data_valid_p9            ( hmc_port[10].wr_data_valid ),
        .hmc_wr_data_ready_p9            ( hmc_port[10].wr_data_ready ),
        .hmc_rd_data_p9                  ( hmc_port[10].rd_data ),
        .hmc_rd_data_tag_p9              ( hmc_port[10].rd_data_tag ),
        .hmc_rd_data_valid_p9            ( hmc_port[10].rd_data_valid ),
        .hmc_errstat_p9                  ( hmc_port[10].errstat ),
        .hmc_dinv_p9                     ( hmc_port[10].dinv ),
        .hmc_clk_p10                     ( hmc_port[11].clk ),
        .hmc_addr_p10                    ( hmc_port[11].addr ),
        .hmc_size_p10                    ( hmc_port[11].size ),
        .hmc_tag_p10                     ( hmc_port[11].tag ),
        .hmc_cmd_valid_p10               ( hmc_port[11].cmd_valid ),
        .hmc_cmd_ready_p10               ( hmc_port[11].cmd_ready ),
        .hmc_cmd_p10                     ( hmc_port[11].cmd ),
        .hmc_wr_data_p10                 ( hmc_port[11].wr_data ),
        .hmc_wr_data_valid_p10           ( hmc_port[11].wr_data_valid ),
        .hmc_wr_data_ready_p10           ( hmc_port[11].wr_data_ready ),
        .hmc_rd_data_p10                 ( hmc_port[11].rd_data ),
        .hmc_rd_data_tag_p10             ( hmc_port[11].rd_data_tag ),
        .hmc_rd_data_valid_p10           ( hmc_port[11].rd_data_valid ),
        .hmc_errstat_p10                 ( hmc_port[11].errstat ),
        .hmc_dinv_p10                    ( hmc_port[11].dinv ),
        .hmc_clk_p11                     ( hmc_port[12].clk ),
        .hmc_addr_p11                    ( hmc_port[12].addr ),
        .hmc_size_p11                    ( hmc_port[12].size ),
        .hmc_tag_p11                     ( hmc_port[12].tag ),
        .hmc_cmd_valid_p11               ( hmc_port[12].cmd_valid ),
        .hmc_cmd_ready_p11               ( hmc_port[12].cmd_ready ),
        .hmc_cmd_p11                     ( hmc_port[12].cmd ),
        .hmc_wr_data_p11                 ( hmc_port[12].wr_data ),
        .hmc_wr_data_valid_p11           ( hmc_port[12].wr_data_valid ),
        .hmc_wr_data_ready_p11           ( hmc_port[12].wr_data_ready ),
        .hmc_rd_data_p11                 ( hmc_port[12].rd_data ),
        .hmc_rd_data_tag_p11             ( hmc_port[12].rd_data_tag ),
        .hmc_rd_data_valid_p11           ( hmc_port[12].rd_data_valid ),
        .hmc_errstat_p11                 ( hmc_port[12].errstat ),
        .hmc_dinv_p11                    ( hmc_port[12].dinv ),
        .hmc_clk_p12                     ( hmc_port[13].clk ),
        .hmc_addr_p12                    ( hmc_port[13].addr ),
        .hmc_size_p12                    ( hmc_port[13].size ),
        .hmc_tag_p12                     ( hmc_port[13].tag ),
        .hmc_cmd_valid_p12               ( hmc_port[13].cmd_valid ),
        .hmc_cmd_ready_p12               ( hmc_port[13].cmd_ready ),
        .hmc_cmd_p12                     ( hmc_port[13].cmd ),
        .hmc_wr_data_p12                 ( hmc_port[13].wr_data ),
        .hmc_wr_data_valid_p12           ( hmc_port[13].wr_data_valid ),
        .hmc_wr_data_ready_p12           ( hmc_port[13].wr_data_ready ),
        .hmc_rd_data_p12                 ( hmc_port[13].rd_data ),
        .hmc_rd_data_tag_p12             ( hmc_port[13].rd_data_tag ),
        .hmc_rd_data_valid_p12           ( hmc_port[13].rd_data_valid ),
        .hmc_errstat_p12                 ( hmc_port[13].errstat ),
        .hmc_dinv_p12                    ( hmc_port[13].dinv ),
        .hmc_clk_p13                     ( hmc_port[14].clk ),
        .hmc_addr_p13                    ( hmc_port[14].addr ),
        .hmc_size_p13                    ( hmc_port[14].size ),
        .hmc_tag_p13                     ( hmc_port[14].tag ),
        .hmc_cmd_valid_p13               ( hmc_port[14].cmd_valid ),
        .hmc_cmd_ready_p13               ( hmc_port[14].cmd_ready ),
        .hmc_cmd_p13                     ( hmc_port[14].cmd ),
        .hmc_wr_data_p13                 ( hmc_port[14].wr_data ),
        .hmc_wr_data_valid_p13           ( hmc_port[14].wr_data_valid ),
        .hmc_wr_data_ready_p13           ( hmc_port[14].wr_data_ready ),
        .hmc_rd_data_p13                 ( hmc_port[14].rd_data ),
        .hmc_rd_data_tag_p13             ( hmc_port[14].rd_data_tag ),
        .hmc_rd_data_valid_p13           ( hmc_port[14].rd_data_valid ),
        .hmc_errstat_p13                 ( hmc_port[14].errstat ),
        .hmc_dinv_p13                    ( hmc_port[14].dinv ),
	  `endif // ENABLE_3RD_HMC_LINK
      `ifdef ENABLE_4TH_HMC_LINK
        .hmc_clk_p14                     ( hmc_port[15].clk ),
        .hmc_addr_p14                    ( hmc_port[15].addr ),
        .hmc_size_p14                    ( hmc_port[15].size ),
        .hmc_tag_p14                     ( hmc_port[15].tag ),
        .hmc_cmd_valid_p14               ( hmc_port[15].cmd_valid ),
        .hmc_cmd_ready_p14               ( hmc_port[15].cmd_ready ),
        .hmc_cmd_p14                     ( hmc_port[15].cmd ),
        .hmc_wr_data_p14                 ( hmc_port[15].wr_data ),
        .hmc_wr_data_valid_p14           ( hmc_port[15].wr_data_valid ),
        .hmc_wr_data_ready_p14           ( hmc_port[15].wr_data_ready ),
        .hmc_rd_data_p14                 ( hmc_port[15].rd_data ),
        .hmc_rd_data_tag_p14             ( hmc_port[15].rd_data_tag ),
        .hmc_rd_data_valid_p14           ( hmc_port[15].rd_data_valid ),
        .hmc_errstat_p14                 ( hmc_port[15].errstat ),
        .hmc_dinv_p14                    ( hmc_port[15].dinv ),
        .hmc_clk_p15                     ( hmc_port[16].clk ),
        .hmc_addr_p15                    ( hmc_port[16].addr ),
        .hmc_size_p15                    ( hmc_port[16].size ),
        .hmc_tag_p15                     ( hmc_port[16].tag ),
        .hmc_cmd_valid_p15               ( hmc_port[16].cmd_valid ),
        .hmc_cmd_ready_p15               ( hmc_port[16].cmd_ready ),
        .hmc_cmd_p15                     ( hmc_port[16].cmd ),
        .hmc_wr_data_p15                 ( hmc_port[16].wr_data ),
        .hmc_wr_data_valid_p15           ( hmc_port[16].wr_data_valid ),
        .hmc_wr_data_ready_p15           ( hmc_port[16].wr_data_ready ),
        .hmc_rd_data_p15                 ( hmc_port[16].rd_data ),
        .hmc_rd_data_tag_p15             ( hmc_port[16].rd_data_tag ),
        .hmc_rd_data_valid_p15           ( hmc_port[16].rd_data_valid ),
        .hmc_errstat_p15                 ( hmc_port[16].errstat ),
        .hmc_dinv_p15                    ( hmc_port[16].dinv ),
        .hmc_clk_p16                     ( hmc_port[17].clk ),
        .hmc_addr_p16                    ( hmc_port[17].addr ),
        .hmc_size_p16                    ( hmc_port[17].size ),
        .hmc_tag_p16                     ( hmc_port[17].tag ),
        .hmc_cmd_valid_p16               ( hmc_port[17].cmd_valid ),
        .hmc_cmd_ready_p16               ( hmc_port[17].cmd_ready ),
        .hmc_cmd_p16                     ( hmc_port[17].cmd ),
        .hmc_wr_data_p16                 ( hmc_port[17].wr_data ),
        .hmc_wr_data_valid_p16           ( hmc_port[17].wr_data_valid ),
        .hmc_wr_data_ready_p16           ( hmc_port[17].wr_data_ready ),
        .hmc_rd_data_p16                 ( hmc_port[17].rd_data ),
        .hmc_rd_data_tag_p16             ( hmc_port[17].rd_data_tag ),
        .hmc_rd_data_valid_p16           ( hmc_port[17].rd_data_valid ),
        .hmc_errstat_p16                 ( hmc_port[17].errstat ),
        .hmc_dinv_p16                    ( hmc_port[17].dinv ),
        .hmc_clk_p17                     ( hmc_port[18].clk ),
        .hmc_addr_p17                    ( hmc_port[18].addr ),
        .hmc_size_p17                    ( hmc_port[18].size ),
        .hmc_tag_p17                     ( hmc_port[18].tag ),
        .hmc_cmd_valid_p17               ( hmc_port[18].cmd_valid ),
        .hmc_cmd_ready_p17               ( hmc_port[18].cmd_ready ),
        .hmc_cmd_p17                     ( hmc_port[18].cmd ),
        .hmc_wr_data_p17                 ( hmc_port[18].wr_data ),
        .hmc_wr_data_valid_p17           ( hmc_port[18].wr_data_valid ),
        .hmc_wr_data_ready_p17           ( hmc_port[18].wr_data_ready ),
        .hmc_rd_data_p17                 ( hmc_port[18].rd_data ),
        .hmc_rd_data_tag_p17             ( hmc_port[18].rd_data_tag ),
        .hmc_rd_data_valid_p17           ( hmc_port[18].rd_data_valid ),
        .hmc_errstat_p17                 ( hmc_port[18].errstat ),
        .hmc_dinv_p17                    ( hmc_port[18].dinv ),
        .hmc_clk_p18                     ( hmc_port[19].clk ),
        .hmc_addr_p18                    ( hmc_port[19].addr ),
        .hmc_size_p18                    ( hmc_port[19].size ),
        .hmc_tag_p18                     ( hmc_port[19].tag ),
        .hmc_cmd_valid_p18               ( hmc_port[19].cmd_valid ),
        .hmc_cmd_ready_p18               ( hmc_port[19].cmd_ready ),
        .hmc_cmd_p18                     ( hmc_port[19].cmd ),
        .hmc_wr_data_p18                 ( hmc_port[19].wr_data ),
        .hmc_wr_data_valid_p18           ( hmc_port[19].wr_data_valid ),
        .hmc_wr_data_ready_p18           ( hmc_port[19].wr_data_ready ),
        .hmc_rd_data_p18                 ( hmc_port[19].rd_data ),
        .hmc_rd_data_tag_p18             ( hmc_port[19].rd_data_tag ),
        .hmc_rd_data_valid_p18           ( hmc_port[19].rd_data_valid ),
        .hmc_errstat_p18                 ( hmc_port[19].errstat ),
        .hmc_dinv_p18                    ( hmc_port[19].dinv ),
	  `endif // ENABLE_4TH_HMC_LINK
    `endif //USE_512_BIT_HMC_CONTROLLER
        .hmc_tx_clk                         (hmc_tx_clk),
        .hmc_rx_clk                         (hmc_rx_clk),
        .hmc_rst                            (hmc_rst),
        .hmc_trained                        (hmc_trained)
`endif // ENABLE_HMC

`ifdef PICO_DDR3_OR_DDR4
        // user multi-port interface
            `ifdef  UM_PREPEND_COMMA , `endif
            `define UM_PREPEND_COMMA

         //---------------------------------------------
         // DDR3 0 AXI

    `ifdef PICO_AXI_PORT_1
         // Slave 1 Interface
         .c0_s1_axi_clk             ( c0_axi_clk    [1] ),

         // Slave Interface Write Address Ports
         .c0_s1_axi_awid            ( c0_axi_awid   [1] ),
         .c0_s1_axi_awaddr          ( c0_axi_awaddr [1] ),
         .c0_s1_axi_awlen           ( c0_axi_awlen  [1] ),
         .c0_s1_axi_awsize          ( c0_axi_awsize [1] ),
         .c0_s1_axi_awburst         ( c0_axi_awburst[1] ),
         .c0_s1_axi_awlock          ( c0_axi_awlock [1] ),
         .c0_s1_axi_awcache         ( c0_axi_awcache[1] ),
         .c0_s1_axi_awprot          ( c0_axi_awprot [1] ),
         .c0_s1_axi_awqos           ( c0_axi_awqos  [1] ),
         .c0_s1_axi_awvalid         ( c0_axi_awvalid[1] ),
         .c0_s1_axi_awready         ( c0_axi_awready[1] ),

         // Slave Interface Write Data Ports
         .c0_s1_axi_wdata           ( c0_axi_wdata  [1] ),
         .c0_s1_axi_wstrb           ( c0_axi_wstrb  [1] ),
         .c0_s1_axi_wlast           ( c0_axi_wlast  [1] ),
         .c0_s1_axi_wvalid          ( c0_axi_wvalid [1] ),
         .c0_s1_axi_wready          ( c0_axi_wready [1] ),

         // Slave Interface Write Response Ports
         .c0_s1_axi_bid             ( c0_axi_bid    [1] ),
         .c0_s1_axi_bresp           ( c0_axi_bresp  [1] ),
         .c0_s1_axi_bvalid          ( c0_axi_bvalid [1] ),
         .c0_s1_axi_bready          ( c0_axi_bready [1] ),

         // Slave Interface Read Address Ports
         .c0_s1_axi_arid            ( c0_axi_arid   [1] ),
         .c0_s1_axi_araddr          ( c0_axi_araddr [1] ),
         .c0_s1_axi_arlen           ( c0_axi_arlen  [1] ),
         .c0_s1_axi_arsize          ( c0_axi_arsize [1] ),
         .c0_s1_axi_arburst         ( c0_axi_arburst[1] ),
         .c0_s1_axi_arlock          ( c0_axi_arlock [1] ),
         .c0_s1_axi_arcache         ( c0_axi_arcache[1] ),
         .c0_s1_axi_arprot          ( c0_axi_arprot [1] ),
         .c0_s1_axi_arqos           ( c0_axi_arqos  [1] ),
         .c0_s1_axi_arvalid         ( c0_axi_arvalid[1] ),
         .c0_s1_axi_arready         ( c0_axi_arready[1] ),

         // Slave Interface Read Data Ports
         .c0_s1_axi_rid             ( c0_axi_rid    [1] ),
         .c0_s1_axi_rdata           ( c0_axi_rdata  [1] ),
         .c0_s1_axi_rresp           ( c0_axi_rresp  [1] ),
         .c0_s1_axi_rlast           ( c0_axi_rlast  [1] ),
         .c0_s1_axi_rvalid          ( c0_axi_rvalid [1] ),
         .c0_s1_axi_rready          ( c0_axi_rready [1] ),
    `endif // PICO_AXI_PORT_1

    `ifdef PICO_AXI_PORT_2
         // Slave 2 Interface
         .c0_s2_axi_clk             ( c0_axi_clk    [2] ),

         // Slave Interface Write Address Ports
         .c0_s2_axi_awid            ( c0_axi_awid   [2] ),
         .c0_s2_axi_awaddr          ( c0_axi_awaddr [2] ),
         .c0_s2_axi_awlen           ( c0_axi_awlen  [2] ),
         .c0_s2_axi_awsize          ( c0_axi_awsize [2] ),
         .c0_s2_axi_awburst         ( c0_axi_awburst[2] ),
         .c0_s2_axi_awlock          ( c0_axi_awlock [2] ),
         .c0_s2_axi_awcache         ( c0_axi_awcache[2] ),
         .c0_s2_axi_awprot          ( c0_axi_awprot [2] ),
         .c0_s2_axi_awqos           ( c0_axi_awqos  [2] ),
         .c0_s2_axi_awvalid         ( c0_axi_awvalid[2] ),
         .c0_s2_axi_awready         ( c0_axi_awready[2] ),

         // Slave Interface Write Data Ports
         .c0_s2_axi_wdata           ( c0_axi_wdata  [2] ),
         .c0_s2_axi_wstrb           ( c0_axi_wstrb  [2] ),
         .c0_s2_axi_wlast           ( c0_axi_wlast  [2] ),
         .c0_s2_axi_wvalid          ( c0_axi_wvalid [2] ),
         .c0_s2_axi_wready          ( c0_axi_wready [2] ),

         // Slave Interface Write Response Ports
         .c0_s2_axi_bid             ( c0_axi_bid    [2] ),
         .c0_s2_axi_bresp           ( c0_axi_bresp  [2] ),
         .c0_s2_axi_bvalid          ( c0_axi_bvalid [2] ),
         .c0_s2_axi_bready          ( c0_axi_bready [2] ),

         // Slave Interface Read Address Ports
         .c0_s2_axi_arid            ( c0_axi_arid   [2] ),
         .c0_s2_axi_araddr          ( c0_axi_araddr [2] ),
         .c0_s2_axi_arlen           ( c0_axi_arlen  [2] ),
         .c0_s2_axi_arsize          ( c0_axi_arsize [2] ),
         .c0_s2_axi_arburst         ( c0_axi_arburst[2] ),
         .c0_s2_axi_arlock          ( c0_axi_arlock [2] ),
         .c0_s2_axi_arcache         ( c0_axi_arcache[2] ),
         .c0_s2_axi_arprot          ( c0_axi_arprot [2] ),
         .c0_s2_axi_arqos           ( c0_axi_arqos  [2] ),
         .c0_s2_axi_arvalid         ( c0_axi_arvalid[2] ),
         .c0_s2_axi_arready         ( c0_axi_arready[2] ),

         // Slave Interface Read Data Ports
         .c0_s2_axi_rid             ( c0_axi_rid    [2] ),
         .c0_s2_axi_rdata           ( c0_axi_rdata  [2] ),
         .c0_s2_axi_rresp           ( c0_axi_rresp  [2] ),
         .c0_s2_axi_rlast           ( c0_axi_rlast  [2] ),
         .c0_s2_axi_rvalid          ( c0_axi_rvalid [2] ),
         .c0_s2_axi_rready          ( c0_axi_rready [2] ),
    `endif // PICO_AXI_PORT_2

    `ifdef PICO_AXI_PORT_3
         // Slave 3 Interface
         .c0_s3_axi_clk             ( c0_axi_clk    [3] ),

         // Slave Interface Write Address Ports
         .c0_s3_axi_awid            ( c0_axi_awid   [3] ),
         .c0_s3_axi_awaddr          ( c0_axi_awaddr [3] ),
         .c0_s3_axi_awlen           ( c0_axi_awlen  [3] ),
         .c0_s3_axi_awsize          ( c0_axi_awsize [3] ),
         .c0_s3_axi_awburst         ( c0_axi_awburst[3] ),
         .c0_s3_axi_awlock          ( c0_axi_awlock [3] ),
         .c0_s3_axi_awcache         ( c0_axi_awcache[3] ),
         .c0_s3_axi_awprot          ( c0_axi_awprot [3] ),
         .c0_s3_axi_awqos           ( c0_axi_awqos  [3] ),
         .c0_s3_axi_awvalid         ( c0_axi_awvalid[3] ),
         .c0_s3_axi_awready         ( c0_axi_awready[3] ),

         // Slave Interface Write Data Ports
         .c0_s3_axi_wdata           ( c0_axi_wdata  [3] ),
         .c0_s3_axi_wstrb           ( c0_axi_wstrb  [3] ),
         .c0_s3_axi_wlast           ( c0_axi_wlast  [3] ),
         .c0_s3_axi_wvalid          ( c0_axi_wvalid [3] ),
         .c0_s3_axi_wready          ( c0_axi_wready [3] ),

         // Slave Interface Write Response Ports
         .c0_s3_axi_bid             ( c0_axi_bid    [3] ),
         .c0_s3_axi_bresp           ( c0_axi_bresp  [3] ),
         .c0_s3_axi_bvalid          ( c0_axi_bvalid [3] ),
         .c0_s3_axi_bready          ( c0_axi_bready [3] ),

         // Slave Interface Read Address Ports
         .c0_s3_axi_arid            ( c0_axi_arid   [3] ),
         .c0_s3_axi_araddr          ( c0_axi_araddr [3] ),
         .c0_s3_axi_arlen           ( c0_axi_arlen  [3] ),
         .c0_s3_axi_arsize          ( c0_axi_arsize [3] ),
         .c0_s3_axi_arburst         ( c0_axi_arburst[3] ),
         .c0_s3_axi_arlock          ( c0_axi_arlock [3] ),
         .c0_s3_axi_arcache         ( c0_axi_arcache[3] ),
         .c0_s3_axi_arprot          ( c0_axi_arprot [3] ),
         .c0_s3_axi_arqos           ( c0_axi_arqos  [3] ),
         .c0_s3_axi_arvalid         ( c0_axi_arvalid[3] ),
         .c0_s3_axi_arready         ( c0_axi_arready[3] ),

         // Slave Interface Read Data Ports
         .c0_s3_axi_rid             ( c0_axi_rid    [3] ),
         .c0_s3_axi_rdata           ( c0_axi_rdata  [3] ),
         .c0_s3_axi_rresp           ( c0_axi_rresp  [3] ),
         .c0_s3_axi_rlast           ( c0_axi_rlast  [3] ),
         .c0_s3_axi_rvalid          ( c0_axi_rvalid [3] ),
         .c0_s3_axi_rready          ( c0_axi_rready [3] ),
    `endif // PICO_AXI_PORT_3

    `ifdef PICO_AXI_PORT_4
         // Slave 4 Interface
         .c0_s4_axi_clk             ( c0_axi_clk    [4] ),

         // Slave Interface Write Address Ports
         .c0_s4_axi_awid            ( c0_axi_awid   [4] ),
         .c0_s4_axi_awaddr          ( c0_axi_awaddr [4] ),
         .c0_s4_axi_awlen           ( c0_axi_awlen  [4] ),
         .c0_s4_axi_awsize          ( c0_axi_awsize [4] ),
         .c0_s4_axi_awburst         ( c0_axi_awburst[4] ),
         .c0_s4_axi_awlock          ( c0_axi_awlock [4] ),
         .c0_s4_axi_awcache         ( c0_axi_awcache[4] ),
         .c0_s4_axi_awprot          ( c0_axi_awprot [4] ),
         .c0_s4_axi_awqos           ( c0_axi_awqos  [4] ),
         .c0_s4_axi_awvalid         ( c0_axi_awvalid[4] ),
         .c0_s4_axi_awready         ( c0_axi_awready[4] ),

         // Slave Interface Write Data Ports
         .c0_s4_axi_wdata           ( c0_axi_wdata  [4] ),
         .c0_s4_axi_wstrb           ( c0_axi_wstrb  [4] ),
         .c0_s4_axi_wlast           ( c0_axi_wlast  [4] ),
         .c0_s4_axi_wvalid          ( c0_axi_wvalid [4] ),
         .c0_s4_axi_wready          ( c0_axi_wready [4] ),

         // Slave Interface Write Response Ports
         .c0_s4_axi_bid             ( c0_axi_bid    [4] ),
         .c0_s4_axi_bresp           ( c0_axi_bresp  [4] ),
         .c0_s4_axi_bvalid          ( c0_axi_bvalid [4] ),
         .c0_s4_axi_bready          ( c0_axi_bready [4] ),

         // Slave Interface Read Address Ports
         .c0_s4_axi_arid            ( c0_axi_arid   [4] ),
         .c0_s4_axi_araddr          ( c0_axi_araddr [4] ),
         .c0_s4_axi_arlen           ( c0_axi_arlen  [4] ),
         .c0_s4_axi_arsize          ( c0_axi_arsize [4] ),
         .c0_s4_axi_arburst         ( c0_axi_arburst[4] ),
         .c0_s4_axi_arlock          ( c0_axi_arlock [4] ),
         .c0_s4_axi_arcache         ( c0_axi_arcache[4] ),
         .c0_s4_axi_arprot          ( c0_axi_arprot [4] ),
         .c0_s4_axi_arqos           ( c0_axi_arqos  [4] ),
         .c0_s4_axi_arvalid         ( c0_axi_arvalid[4] ),
         .c0_s4_axi_arready         ( c0_axi_arready[4] ),

         // Slave Interface Read Data Ports
         .c0_s4_axi_rid             ( c0_axi_rid    [4] ),
         .c0_s4_axi_rdata           ( c0_axi_rdata  [4] ),
         .c0_s4_axi_rresp           ( c0_axi_rresp  [4] ),
         .c0_s4_axi_rlast           ( c0_axi_rlast  [4] ),
         .c0_s4_axi_rvalid          ( c0_axi_rvalid [4] ),
         .c0_s4_axi_rready          ( c0_axi_rready [4] ),
    `endif // PICO_AXI_PORT_4

    `ifdef PICO_AXI_PORT_5
         // Slave 5 Interface
         .c0_s5_axi_clk             ( c0_axi_clk    [5] ),

         // Slave Interface Write Address Ports
         .c0_s5_axi_awid            ( c0_axi_awid   [5] ),
         .c0_s5_axi_awaddr          ( c0_axi_awaddr [5] ),
         .c0_s5_axi_awlen           ( c0_axi_awlen  [5] ),
         .c0_s5_axi_awsize          ( c0_axi_awsize [5] ),
         .c0_s5_axi_awburst         ( c0_axi_awburst[5] ),
         .c0_s5_axi_awlock          ( c0_axi_awlock [5] ),
         .c0_s5_axi_awcache         ( c0_axi_awcache[5] ),
         .c0_s5_axi_awprot          ( c0_axi_awprot [5] ),
         .c0_s5_axi_awqos           ( c0_axi_awqos  [5] ),
         .c0_s5_axi_awvalid         ( c0_axi_awvalid[5] ),
         .c0_s5_axi_awready         ( c0_axi_awready[5] ),

         // Slave Interface Write Data Ports
         .c0_s5_axi_wdata           ( c0_axi_wdata  [5] ),
         .c0_s5_axi_wstrb           ( c0_axi_wstrb  [5] ),
         .c0_s5_axi_wlast           ( c0_axi_wlast  [5] ),
         .c0_s5_axi_wvalid          ( c0_axi_wvalid [5] ),
         .c0_s5_axi_wready          ( c0_axi_wready [5] ),

         // Slave Interface Write Response Ports
         .c0_s5_axi_bid             ( c0_axi_bid    [5] ),
         .c0_s5_axi_bresp           ( c0_axi_bresp  [5] ),
         .c0_s5_axi_bvalid          ( c0_axi_bvalid [5] ),
         .c0_s5_axi_bready          ( c0_axi_bready [5] ),

         // Slave Interface Read Address Ports
         .c0_s5_axi_arid            ( c0_axi_arid   [5] ),
         .c0_s5_axi_araddr          ( c0_axi_araddr [5] ),
         .c0_s5_axi_arlen           ( c0_axi_arlen  [5] ),
         .c0_s5_axi_arsize          ( c0_axi_arsize [5] ),
         .c0_s5_axi_arburst         ( c0_axi_arburst[5] ),
         .c0_s5_axi_arlock          ( c0_axi_arlock [5] ),
         .c0_s5_axi_arcache         ( c0_axi_arcache[5] ),
         .c0_s5_axi_arprot          ( c0_axi_arprot [5] ),
         .c0_s5_axi_arqos           ( c0_axi_arqos  [5] ),
         .c0_s5_axi_arvalid         ( c0_axi_arvalid[5] ),
         .c0_s5_axi_arready         ( c0_axi_arready[5] ),

         // Slave Interface Read Data Ports
         .c0_s5_axi_rid             ( c0_axi_rid    [5] ),
         .c0_s5_axi_rdata           ( c0_axi_rdata  [5] ),
         .c0_s5_axi_rresp           ( c0_axi_rresp  [5] ),
         .c0_s5_axi_rlast           ( c0_axi_rlast  [5] ),
         .c0_s5_axi_rvalid          ( c0_axi_rvalid [5] ),
         .c0_s5_axi_rready          ( c0_axi_rready [5] ),
    `endif // PICO_AXI_PORT_5

    `ifdef PICO_AXI_PORT_6
         // Slave 6 Interface
         .c0_s6_axi_clk             ( c0_axi_clk    [6] ),

         // Slave Interface Write Address Ports
         .c0_s6_axi_awid            ( c0_axi_awid   [6] ),
         .c0_s6_axi_awaddr          ( c0_axi_awaddr [6] ),
         .c0_s6_axi_awlen           ( c0_axi_awlen  [6] ),
         .c0_s6_axi_awsize          ( c0_axi_awsize [6] ),
         .c0_s6_axi_awburst         ( c0_axi_awburst[6] ),
         .c0_s6_axi_awlock          ( c0_axi_awlock [6] ),
         .c0_s6_axi_awcache         ( c0_axi_awcache[6] ),
         .c0_s6_axi_awprot          ( c0_axi_awprot [6] ),
         .c0_s6_axi_awqos           ( c0_axi_awqos  [6] ),
         .c0_s6_axi_awvalid         ( c0_axi_awvalid[6] ),
         .c0_s6_axi_awready         ( c0_axi_awready[6] ),

         // Slave Interface Write Data Ports
         .c0_s6_axi_wdata           ( c0_axi_wdata  [6] ),
         .c0_s6_axi_wstrb           ( c0_axi_wstrb  [6] ),
         .c0_s6_axi_wlast           ( c0_axi_wlast  [6] ),
         .c0_s6_axi_wvalid          ( c0_axi_wvalid [6] ),
         .c0_s6_axi_wready          ( c0_axi_wready [6] ),

         // Slave Interface Write Response Ports
         .c0_s6_axi_bid             ( c0_axi_bid    [6] ),
         .c0_s6_axi_bresp           ( c0_axi_bresp  [6] ),
         .c0_s6_axi_bvalid          ( c0_axi_bvalid [6] ),
         .c0_s6_axi_bready          ( c0_axi_bready [6] ),

         // Slave Interface Read Address Ports
         .c0_s6_axi_arid            ( c0_axi_arid   [6] ),
         .c0_s6_axi_araddr          ( c0_axi_araddr [6] ),
         .c0_s6_axi_arlen           ( c0_axi_arlen  [6] ),
         .c0_s6_axi_arsize          ( c0_axi_arsize [6] ),
         .c0_s6_axi_arburst         ( c0_axi_arburst[6] ),
         .c0_s6_axi_arlock          ( c0_axi_arlock [6] ),
         .c0_s6_axi_arcache         ( c0_axi_arcache[6] ),
         .c0_s6_axi_arprot          ( c0_axi_arprot [6] ),
         .c0_s6_axi_arqos           ( c0_axi_arqos  [6] ),
         .c0_s6_axi_arvalid         ( c0_axi_arvalid[6] ),
         .c0_s6_axi_arready         ( c0_axi_arready[6] ),

         // Slave Interface Read Data Ports
         .c0_s6_axi_rid             ( c0_axi_rid    [6] ),
         .c0_s6_axi_rdata           ( c0_axi_rdata  [6] ),
         .c0_s6_axi_rresp           ( c0_axi_rresp  [6] ),
         .c0_s6_axi_rlast           ( c0_axi_rlast  [6] ),
         .c0_s6_axi_rvalid          ( c0_axi_rvalid [6] ),
         .c0_s6_axi_rready          ( c0_axi_rready [6] ),
    `endif // PICO_AXI_PORT_6

    `ifdef PICO_AXI_PORT_7
         // Slave 7 Interface
         .c0_s7_axi_clk             ( c0_axi_clk    [7] ),

         // Slave Interface Write Address Ports
         .c0_s7_axi_awid            ( c0_axi_awid   [7] ),
         .c0_s7_axi_awaddr          ( c0_axi_awaddr [7] ),
         .c0_s7_axi_awlen           ( c0_axi_awlen  [7] ),
         .c0_s7_axi_awsize          ( c0_axi_awsize [7] ),
         .c0_s7_axi_awburst         ( c0_axi_awburst[7] ),
         .c0_s7_axi_awlock          ( c0_axi_awlock [7] ),
         .c0_s7_axi_awcache         ( c0_axi_awcache[7] ),
         .c0_s7_axi_awprot          ( c0_axi_awprot [7] ),
         .c0_s7_axi_awqos           ( c0_axi_awqos  [7] ),
         .c0_s7_axi_awvalid         ( c0_axi_awvalid[7] ),
         .c0_s7_axi_awready         ( c0_axi_awready[7] ),

         // Slave Interface Write Data Ports
         .c0_s7_axi_wdata           ( c0_axi_wdata  [7] ),
         .c0_s7_axi_wstrb           ( c0_axi_wstrb  [7] ),
         .c0_s7_axi_wlast           ( c0_axi_wlast  [7] ),
         .c0_s7_axi_wvalid          ( c0_axi_wvalid [7] ),
         .c0_s7_axi_wready          ( c0_axi_wready [7] ),

         // Slave Interface Write Response Ports
         .c0_s7_axi_bid             ( c0_axi_bid    [7] ),
         .c0_s7_axi_bresp           ( c0_axi_bresp  [7] ),
         .c0_s7_axi_bvalid          ( c0_axi_bvalid [7] ),
         .c0_s7_axi_bready          ( c0_axi_bready [7] ),

         // Slave Interface Read Address Ports
         .c0_s7_axi_arid            ( c0_axi_arid   [7] ),
         .c0_s7_axi_araddr          ( c0_axi_araddr [7] ),
         .c0_s7_axi_arlen           ( c0_axi_arlen  [7] ),
         .c0_s7_axi_arsize          ( c0_axi_arsize [7] ),
         .c0_s7_axi_arburst         ( c0_axi_arburst[7] ),
         .c0_s7_axi_arlock          ( c0_axi_arlock [7] ),
         .c0_s7_axi_arcache         ( c0_axi_arcache[7] ),
         .c0_s7_axi_arprot          ( c0_axi_arprot [7] ),
         .c0_s7_axi_arqos           ( c0_axi_arqos  [7] ),
         .c0_s7_axi_arvalid         ( c0_axi_arvalid[7] ),
         .c0_s7_axi_arready         ( c0_axi_arready[7] ),

         // Slave Interface Read Data Ports
         .c0_s7_axi_rid             ( c0_axi_rid    [7] ),
         .c0_s7_axi_rdata           ( c0_axi_rdata  [7] ),
         .c0_s7_axi_rresp           ( c0_axi_rresp  [7] ),
         .c0_s7_axi_rlast           ( c0_axi_rlast  [7] ),
         .c0_s7_axi_rvalid          ( c0_axi_rvalid [7] ),
         .c0_s7_axi_rready          ( c0_axi_rready [7] ),
    `endif // PICO_AXI_PORT_7

         // AXI clock and reset
         `ifndef PICO_MODEL_SB852
         .c0_axi_clk                ( c0_tb_clk         ),
         .c0_axi_rst                ( c0_tb_rst         ),
         `else
         .c0_axi_clk                ( c0_clk            ),
         .c0_axi_rst                ( c0_rst            ),
         `endif
         .c0_phy_init_done          ( c0_phy_init_done  )
`endif //PICO_DDR3_OR_DDR4

    // Below are ifdefs with the stream signals being brought in.
    // Copy the names from the stream1 and change the 1 to what you are bringing in, format is the same throughout
    `ifdef STREAM1_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s1i_rdy(stream_in_rdy[1]),
        .s1i_valid(stream_in_valid[1]),
    `ifdef STREAM1_IN_256BIT
	.s1i_ow_dvld(stream_in_ow_dvld[1][OW_DVLD_W-1:0]),
    `endif
        .s1i_data(stream_in_data[1][`STREAM1_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM1_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s1o_rdy(stream_out_rdy[1]),
        .s1o_valid(stream_out_valid[1]),
    `ifdef STREAM1_OUT_256BIT
	.s1o_ow_dvld(stream_out_ow_dvld[1][OW_DVLD_W-1:0]),
    `endif
        .s1o_data(stream_out_data[1][`STREAM1_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM2_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s2i_rdy(stream_in_rdy[2]),
        .s2i_valid(stream_in_valid[2]),
    `ifdef STREAM2_IN_256BIT
	.s2i_ow_dvld(stream_in_ow_dvld[2][OW_DVLD_W-1:0]),
    `endif
        .s2i_data(stream_in_data[2][`STREAM2_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM2_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s2o_rdy(stream_out_rdy[2]),
        .s2o_valid(stream_out_valid[2]),
    `ifdef STREAM2_OUT_256BIT
	.s2o_ow_dvld(stream_out_ow_dvld[2][OW_DVLD_W-1:0]),
    `endif
        .s2o_data(stream_out_data[2][`STREAM2_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM3_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s3i_rdy(stream_in_rdy[3]),
        .s3i_valid(stream_in_valid[3]),
    `ifdef STREAM3_IN_256BIT
	.s3i_ow_dvld(stream_in_ow_dvld[3][OW_DVLD_W-1:0]),
    `endif
        .s3i_data(stream_in_data[3][`STREAM3_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM3_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s3o_rdy(stream_out_rdy[3]),
        .s3o_valid(stream_out_valid[3]),
    `ifdef STREAM3_OUT_256BIT
	.s3o_ow_dvld(stream_out_ow_dvld[3][OW_DVLD_W-1:0]),
    `endif
        .s3o_data(stream_out_data[3][`STREAM3_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM4_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s4i_rdy(stream_in_rdy[4]),
        .s4i_valid(stream_in_valid[4]),
    `ifdef STREAM4_IN_256BIT
	.s4i_ow_dvld(stream_in_ow_dvld[4][OW_DVLD_W-1:0]),
    `endif
        .s4i_data(stream_in_data[4][`STREAM4_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM4_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s4o_rdy(stream_out_rdy[4]),
        .s4o_valid(stream_out_valid[4]),
    `ifdef STREAM4_OUT_256BIT
	.s4o_ow_dvld(stream_out_ow_dvld[4][OW_DVLD_W-1:0]),
    `endif
        .s4o_data(stream_out_data[4][`STREAM4_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM5_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s5i_rdy(stream_in_rdy[5]),
        .s5i_valid(stream_in_valid[5]),
    `ifdef STREAM5_IN_256BIT
	.s5i_ow_dvld(stream_in_ow_dvld[5][OW_DVLD_W-1:0]),
    `endif
        .s5i_data(stream_in_data[5][`STREAM5_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM5_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s5o_rdy(stream_out_rdy[5]),
        .s5o_valid(stream_out_valid[5]),
    `ifdef STREAM5_OUT_256BIT
	.s5o_ow_dvld(stream_out_ow_dvld[5][OW_DVLD_W-1:0]),
    `endif
        .s5o_data(stream_out_data[5][`STREAM5_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM6_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s6i_rdy(stream_in_rdy[6]),
        .s6i_valid(stream_in_valid[6]),
    `ifdef STREAM6_IN_256BIT
	.s6i_ow_dvld(stream_in_ow_dvld[6][OW_DVLD_W-1:0]),
    `endif
        .s6i_data(stream_in_data[6][`STREAM6_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM6_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s6o_rdy(stream_out_rdy[6]),
        .s6o_valid(stream_out_valid[6]),
    `ifdef STREAM6_OUT_256BIT
	.s6o_ow_dvld(stream_out_ow_dvld[6][OW_DVLD_W-1:0]),
    `endif
        .s6o_data(stream_out_data[6][`STREAM6_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM7_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s7i_rdy(stream_in_rdy[7]),
        .s7i_valid(stream_in_valid[7]),
    `ifdef STREAM7_IN_256BIT
	.s7i_ow_dvld(stream_in_ow_dvld[7][OW_DVLD_W-1:0]),
    `endif
        .s7i_data(stream_in_data[7][`STREAM7_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM7_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s7o_rdy(stream_out_rdy[7]),
        .s7o_valid(stream_out_valid[7]),
    `ifdef STREAM7_OUT_256BIT
	.s7o_ow_dvld(stream_out_ow_dvld[7][OW_DVLD_W-1:0]),
    `endif
        .s7o_data(stream_out_data[7][`STREAM7_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM8_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s8i_rdy(stream_in_rdy[8]),
        .s8i_valid(stream_in_valid[8]),
    `ifdef STREAM8_IN_256BIT
	.s8i_ow_dvld(stream_in_ow_dvld[8][OW_DVLD_W-1:0]),
    `endif
        .s8i_data(stream_in_data[8][`STREAM8_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM8_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s8o_rdy(stream_out_rdy[8]),
        .s8o_valid(stream_out_valid[8]),
    `ifdef STREAM8_OUT_256BIT
	.s8o_ow_dvld(stream_out_ow_dvld[8][OW_DVLD_W-1:0]),
    `endif
        .s8o_data(stream_out_data[8][`STREAM8_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM9_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s9i_rdy(stream_in_rdy[9]),
        .s9i_valid(stream_in_valid[9]),
    `ifdef STREAM9_IN_256BIT
	.s9i_ow_dvld(stream_in_ow_dvld[9][OW_DVLD_W-1:0]),
    `endif
        .s9i_data(stream_in_data[9][`STREAM9_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM9_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s9o_rdy(stream_out_rdy[9]),
        .s9o_valid(stream_out_valid[9]),
    `ifdef STREAM9_OUT_256BIT
	.s9o_ow_dvld(stream_out_ow_dvld[9][OW_DVLD_W-1:0]),
    `endif
        .s9o_data(stream_out_data[9][`STREAM9_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM10_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s10i_rdy(stream_in_rdy[10]),
        .s10i_valid(stream_in_valid[10]),
    `ifdef STREAM10_IN_256BIT
	.s10i_ow_dvld(stream_in_ow_dvld[10][OW_DVLD_W-1:0]),
    `endif
        .s10i_data(stream_in_data[10][`STREAM10_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM10_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s10o_rdy(stream_out_rdy[10]),
        .s10o_valid(stream_out_valid[10]),
    `ifdef STREAM10_OUT_256BIT
	.s10o_ow_dvld(stream_out_ow_dvld[10][OW_DVLD_W-1:0]),
    `endif
        .s10o_data(stream_out_data[10][`STREAM10_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM11_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s11i_rdy(stream_in_rdy[11]),
        .s11i_valid(stream_in_valid[11]),
    `ifdef STREAM11_IN_256BIT
	.s11i_ow_dvld(stream_in_ow_dvld[11][OW_DVLD_W-1:0]),
    `endif
        .s11i_data(stream_in_data[11][`STREAM11_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM11_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s11o_rdy(stream_out_rdy[11]),
        .s11o_valid(stream_out_valid[11]),
    `ifdef STREAM11_OUT_256BIT
	.s11o_ow_dvld(stream_out_ow_dvld[11][OW_DVLD_W-1:0]),
    `endif
        .s11o_data(stream_out_data[11][`STREAM11_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM12_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s12i_rdy(stream_in_rdy[12]),
        .s12i_valid(stream_in_valid[12]),
    `ifdef STREAM12_IN_256BIT
	.s12i_ow_dvld(stream_in_ow_dvld[12][OW_DVLD_W-1:0]),
    `endif
        .s12i_data(stream_in_data[12][`STREAM12_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM12_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s12o_rdy(stream_out_rdy[12]),
        .s12o_valid(stream_out_valid[12]),
    `ifdef STREAM12_OUT_256BIT
	.s12o_ow_dvld(stream_out_ow_dvld[12][OW_DVLD_W-1:0]),
    `endif
        .s12o_data(stream_out_data[12][`STREAM12_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM13_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s13i_rdy(stream_in_rdy[13]),
        .s13i_valid(stream_in_valid[13]),
    `ifdef STREAM13_IN_256BIT
	.s13i_ow_dvld(stream_in_ow_dvld[13][OW_DVLD_W-1:0]),
    `endif
        .s13i_data(stream_in_data[13][`STREAM13_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM13_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s13o_rdy(stream_out_rdy[13]),
        .s13o_valid(stream_out_valid[13]),
    `ifdef STREAM13_OUT_256BIT
	.s13o_ow_dvld(stream_out_ow_dvld[13][OW_DVLD_W-1:0]),
    `endif
        .s13o_data(stream_out_data[13][`STREAM13_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM14_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s14i_rdy(stream_in_rdy[14]),
        .s14i_valid(stream_in_valid[14]),
    `ifdef STREAM14_IN_256BIT
	.s14i_ow_dvld(stream_in_ow_dvld[14][OW_DVLD_W-1:0]),
    `endif
        .s14i_data(stream_in_data[14][`STREAM14_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM14_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s14o_rdy(stream_out_rdy[14]),
        .s14o_valid(stream_out_valid[14]),
    `ifdef STREAM14_OUT_256BIT
	.s14o_ow_dvld(stream_out_ow_dvld[14][OW_DVLD_W-1:0]),
    `endif
        .s14o_data(stream_out_data[14][`STREAM14_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM15_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s15i_rdy(stream_in_rdy[15]),
        .s15i_valid(stream_in_valid[15]),
    `ifdef STREAM15_IN_256BIT
	.s15i_ow_dvld(stream_in_ow_dvld[15][OW_DVLD_W-1:0]),
    `endif
        .s15i_data(stream_in_data[15][`STREAM15_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM15_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s15o_rdy(stream_out_rdy[15]),
        .s15o_valid(stream_out_valid[15]),
    `ifdef STREAM15_OUT_256BIT
	.s15o_ow_dvld(stream_out_ow_dvld[15][OW_DVLD_W-1:0]),
    `endif
        .s15o_data(stream_out_data[15][`STREAM15_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM16_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s16i_rdy(stream_in_rdy[16]),
        .s16i_valid(stream_in_valid[16]),
    `ifdef STREAM16_IN_256BIT
	.s16i_ow_dvld(stream_in_ow_dvld[16][OW_DVLD_W-1:0]),
    `endif
        .s16i_data(stream_in_data[16][`STREAM16_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM16_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s16o_rdy(stream_out_rdy[16]),
        .s16o_valid(stream_out_valid[16]),
    `ifdef STREAM16_OUT_256BIT
	.s16o_ow_dvld(stream_out_ow_dvld[16][OW_DVLD_W-1:0]),
    `endif
        .s16o_data(stream_out_data[16][`STREAM16_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM17_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s17i_rdy(stream_in_rdy[17]),
        .s17i_valid(stream_in_valid[17]),
    `ifdef STREAM17_IN_256BIT
	.s17i_ow_dvld(stream_in_ow_dvld[17][OW_DVLD_W-1:0]),
    `endif
        .s17i_data(stream_in_data[17][`STREAM17_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM17_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s17o_rdy(stream_out_rdy[17]),
        .s17o_valid(stream_out_valid[17]),
    `ifdef STREAM17_OUT_256BIT
	.s17o_ow_dvld(stream_out_ow_dvld[17][OW_DVLD_W-1:0]),
    `endif
        .s17o_data(stream_out_data[17][`STREAM17_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM18_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s18i_rdy(stream_in_rdy[18]),
        .s18i_valid(stream_in_valid[18]),
    `ifdef STREAM18_IN_256BIT
	.s18i_ow_dvld(stream_in_ow_dvld[18][OW_DVLD_W-1:0]),
    `endif
        .s18i_data(stream_in_data[18][`STREAM18_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM18_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s18o_rdy(stream_out_rdy[18]),
        .s18o_valid(stream_out_valid[18]),
    `ifdef STREAM18_OUT_256BIT
	.s18o_ow_dvld(stream_out_ow_dvld[18][OW_DVLD_W-1:0]),
    `endif
        .s18o_data(stream_out_data[18][`STREAM18_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM19_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s19i_rdy(stream_in_rdy[19]),
        .s19i_valid(stream_in_valid[19]),
    `ifdef STREAM19_IN_256BIT
	.s19i_ow_dvld(stream_in_ow_dvld[19][OW_DVLD_W-1:0]),
    `endif
        .s19i_data(stream_in_data[19][`STREAM19_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM19_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s19o_rdy(stream_out_rdy[19]),
        .s19o_valid(stream_out_valid[19]),
    `ifdef STREAM19_OUT_256BIT
	.s19o_ow_dvld(stream_out_ow_dvld[19][OW_DVLD_W-1:0]),
    `endif
        .s19o_data(stream_out_data[19][`STREAM19_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM20_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s20i_rdy(stream_in_rdy[20]),
        .s20i_valid(stream_in_valid[20]),
    `ifdef STREAM20_IN_256BIT
	.s20i_ow_dvld(stream_in_ow_dvld[20][OW_DVLD_W-1:0]),
    `endif
        .s20i_data(stream_in_data[20][`STREAM20_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM20_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s20o_rdy(stream_out_rdy[20]),
        .s20o_valid(stream_out_valid[20]),
    `ifdef STREAM20_OUT_256BIT
	.s20o_ow_dvld(stream_out_ow_dvld[20][OW_DVLD_W-1:0]),
    `endif
        .s20o_data(stream_out_data[20][`STREAM20_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM21_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s21i_rdy(stream_in_rdy[21]),
        .s21i_valid(stream_in_valid[21]),
    `ifdef STREAM21_IN_256BIT
	.s21i_ow_dvld(stream_in_ow_dvld[21][OW_DVLD_W-1:0]),
    `endif
        .s21i_data(stream_in_data[21][`STREAM21_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM21_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s21o_rdy(stream_out_rdy[21]),
        .s21o_valid(stream_out_valid[21]),
    `ifdef STREAM21_OUT_256BIT
	.s21o_ow_dvld(stream_out_ow_dvld[21][OW_DVLD_W-1:0]),
    `endif
        .s21o_data(stream_out_data[21][`STREAM21_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM22_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s22i_rdy(stream_in_rdy[22]),
        .s22i_valid(stream_in_valid[22]),
    `ifdef STREAM22_IN_256BIT
	.s22i_ow_dvld(stream_in_ow_dvld[22][OW_DVLD_W-1:0]),
    `endif
        .s22i_data(stream_in_data[22][`STREAM22_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM22_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s22o_rdy(stream_out_rdy[22]),
        .s22o_valid(stream_out_valid[22]),
    `ifdef STREAM22_OUT_256BIT
	.s22o_ow_dvld(stream_out_ow_dvld[22][OW_DVLD_W-1:0]),
    `endif
        .s22o_data(stream_out_data[22][`STREAM22_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM23_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s23i_rdy(stream_in_rdy[23]),
        .s23i_valid(stream_in_valid[23]),
    `ifdef STREAM23_IN_256BIT
	.s23i_ow_dvld(stream_in_ow_dvld[23][OW_DVLD_W-1:0]),
    `endif
        .s23i_data(stream_in_data[23][`STREAM23_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM23_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s23o_rdy(stream_out_rdy[23]),
        .s23o_valid(stream_out_valid[23]),
    `ifdef STREAM23_OUT_256BIT
	.s23o_ow_dvld(stream_out_ow_dvld[23][OW_DVLD_W-1:0]),
    `endif
        .s23o_data(stream_out_data[23][`STREAM23_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM24_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s24i_rdy(stream_in_rdy[24]),
        .s24i_valid(stream_in_valid[24]),
    `ifdef STREAM24_IN_256BIT
	.s24i_ow_dvld(stream_in_ow_dvld[24][OW_DVLD_W-1:0]),
    `endif
        .s24i_data(stream_in_data[24][`STREAM24_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM24_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s24o_rdy(stream_out_rdy[24]),
        .s24o_valid(stream_out_valid[24]),
    `ifdef STREAM24_OUT_256BIT
	.s24o_ow_dvld(stream_out_ow_dvld[24][OW_DVLD_W-1:0]),
    `endif
        .s24o_data(stream_out_data[24][`STREAM24_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM25_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s25i_rdy(stream_in_rdy[25]),
        .s25i_valid(stream_in_valid[25]),
    `ifdef STREAM25_IN_256BIT
	.s25i_ow_dvld(stream_in_ow_dvld[25][OW_DVLD_W-1:0]),
    `endif
        .s25i_data(stream_in_data[25][`STREAM25_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM25_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s25o_rdy(stream_out_rdy[25]),
        .s25o_valid(stream_out_valid[25]),
    `ifdef STREAM25_OUT_256BIT
	.s25o_ow_dvld(stream_out_ow_dvld[25][OW_DVLD_W-1:0]),
    `endif
        .s25o_data(stream_out_data[25][`STREAM25_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM26_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s26i_rdy(stream_in_rdy[26]),
        .s26i_valid(stream_in_valid[26]),
    `ifdef STREAM26_IN_256BIT
	.s26i_ow_dvld(stream_in_ow_dvld[26][OW_DVLD_W-1:0]),
    `endif
        .s26i_data(stream_in_data[26][`STREAM26_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM26_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s26o_rdy(stream_out_rdy[26]),
        .s26o_valid(stream_out_valid[26]),
    `ifdef STREAM26_OUT_256BIT
	.s26o_ow_dvld(stream_out_ow_dvld[26][OW_DVLD_W-1:0]),
    `endif
        .s26o_data(stream_out_data[26][`STREAM26_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM27_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s27i_rdy(stream_in_rdy[27]),
        .s27i_valid(stream_in_valid[27]),
    `ifdef STREAM27_IN_256BIT
	.s27i_ow_dvld(stream_in_ow_dvld[27][OW_DVLD_W-1:0]),
    `endif
        .s27i_data(stream_in_data[27][`STREAM27_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM27_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s27o_rdy(stream_out_rdy[27]),
        .s27o_valid(stream_out_valid[27]),
    `ifdef STREAM27_OUT_256BIT
	.s27o_ow_dvld(stream_out_ow_dvld[27][OW_DVLD_W-1:0]),
    `endif
        .s27o_data(stream_out_data[27][`STREAM27_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM28_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s28i_rdy(stream_in_rdy[28]),
        .s28i_valid(stream_in_valid[28]),
    `ifdef STREAM28_IN_256BIT
	.s28i_ow_dvld(stream_in_ow_dvld[28][OW_DVLD_W-1:0]),
    `endif
        .s28i_data(stream_in_data[28][`STREAM28_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM28_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s28o_rdy(stream_out_rdy[28]),
        .s28o_valid(stream_out_valid[28]),
    `ifdef STREAM28_OUT_256BIT
	.s28o_ow_dvld(stream_out_ow_dvld[28][OW_DVLD_W-1:0]),
    `endif
        .s28o_data(stream_out_data[28][`STREAM28_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM29_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s29i_rdy(stream_in_rdy[29]),
        .s29i_valid(stream_in_valid[29]),
    `ifdef STREAM29_IN_256BIT
	.s29i_ow_dvld(stream_in_ow_dvld[29][OW_DVLD_W-1:0]),
    `endif
        .s29i_data(stream_in_data[29][`STREAM29_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM29_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s29o_rdy(stream_out_rdy[29]),
        .s29o_valid(stream_out_valid[29]),
    `ifdef STREAM29_OUT_256BIT
	.s29o_ow_dvld(stream_out_ow_dvld[29][OW_DVLD_W-1:0]),
    `endif
        .s29o_data(stream_out_data[29][`STREAM29_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM30_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s30i_rdy(stream_in_rdy[30]),
        .s30i_valid(stream_in_valid[30]),
    `ifdef STREAM30_IN_256BIT
	.s30i_ow_dvld(stream_in_ow_dvld[30][OW_DVLD_W-1:0]),
    `endif
        .s30i_data(stream_in_data[30][`STREAM30_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM30_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s30o_rdy(stream_out_rdy[30]),
        .s30o_valid(stream_out_valid[30]),
    `ifdef STREAM30_OUT_256BIT
	.s30o_ow_dvld(stream_out_ow_dvld[30][OW_DVLD_W-1:0]),
    `endif
        .s30o_data(stream_out_data[30][`STREAM30_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM31_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s31i_rdy(stream_in_rdy[31]),
        .s31i_valid(stream_in_valid[31]),
    `ifdef STREAM31_IN_256BIT
	.s31i_ow_dvld(stream_in_ow_dvld[31][OW_DVLD_W-1:0]),
    `endif
        .s31i_data(stream_in_data[31][`STREAM31_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM31_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s31o_rdy(stream_out_rdy[31]),
        .s31o_valid(stream_out_valid[31]),
    `ifdef STREAM31_OUT_256BIT
	.s31o_ow_dvld(stream_out_ow_dvld[31][OW_DVLD_W-1:0]),
    `endif
        .s31o_data(stream_out_data[31][`STREAM31_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM32_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s32i_rdy(stream_in_rdy[32]),
        .s32i_valid(stream_in_valid[32]),
    `ifdef STREAM32_IN_256BIT
	.s32i_ow_dvld(stream_in_ow_dvld[32][OW_DVLD_W-1:0]),
    `endif
        .s32i_data(stream_in_data[32][`STREAM32_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM32_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s32o_rdy(stream_out_rdy[32]),
        .s32o_valid(stream_out_valid[32]),
    `ifdef STREAM32_OUT_256BIT
	.s32o_ow_dvld(stream_out_ow_dvld[32][OW_DVLD_W-1:0]),
    `endif
        .s32o_data(stream_out_data[32][`STREAM32_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM33_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s33i_rdy(stream_in_rdy[33]),
        .s33i_valid(stream_in_valid[33]),
    `ifdef STREAM33_IN_256BIT
	.s33i_ow_dvld(stream_in_ow_dvld[33][OW_DVLD_W-1:0]),
    `endif
        .s33i_data(stream_in_data[33][`STREAM33_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM33_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s33o_rdy(stream_out_rdy[33]),
        .s33o_valid(stream_out_valid[33]),
    `ifdef STREAM33_OUT_256BIT
	.s33o_ow_dvld(stream_out_ow_dvld[33][OW_DVLD_W-1:0]),
    `endif
        .s33o_data(stream_out_data[33][`STREAM33_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM34_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s34i_rdy(stream_in_rdy[34]),
        .s34i_valid(stream_in_valid[34]),
    `ifdef STREAM34_IN_256BIT
	.s34i_ow_dvld(stream_in_ow_dvld[34][OW_DVLD_W-1:0]),
    `endif
        .s34i_data(stream_in_data[34][`STREAM34_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM34_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s34o_rdy(stream_out_rdy[34]),
        .s34o_valid(stream_out_valid[34]),
    `ifdef STREAM34_OUT_256BIT
	.s34o_ow_dvld(stream_out_ow_dvld[34][OW_DVLD_W-1:0]),
    `endif
        .s34o_data(stream_out_data[34][`STREAM34_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM35_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s35i_rdy(stream_in_rdy[35]),
        .s35i_valid(stream_in_valid[35]),
    `ifdef STREAM35_IN_256BIT
	.s35i_ow_dvld(stream_in_ow_dvld[35][OW_DVLD_W-1:0]),
    `endif
        .s35i_data(stream_in_data[35][`STREAM35_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM35_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s35o_rdy(stream_out_rdy[35]),
        .s35o_valid(stream_out_valid[35]),
    `ifdef STREAM35_OUT_256BIT
	.s35o_ow_dvld(stream_out_ow_dvld[35][OW_DVLD_W-1:0]),
    `endif
        .s35o_data(stream_out_data[35][`STREAM35_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM36_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s36i_rdy(stream_in_rdy[36]),
        .s36i_valid(stream_in_valid[36]),
    `ifdef STREAM36_IN_256BIT
	.s36i_ow_dvld(stream_in_ow_dvld[36][OW_DVLD_W-1:0]),
    `endif
        .s36i_data(stream_in_data[36][`STREAM36_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM36_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s36o_rdy(stream_out_rdy[36]),
        .s36o_valid(stream_out_valid[36]),
    `ifdef STREAM36_OUT_256BIT
	.s36o_ow_dvld(stream_out_ow_dvld[36][OW_DVLD_W-1:0]),
    `endif
        .s36o_data(stream_out_data[36][`STREAM36_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM37_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s37i_rdy(stream_in_rdy[37]),
        .s37i_valid(stream_in_valid[37]),
    `ifdef STREAM37_IN_256BIT
	.s37i_ow_dvld(stream_in_ow_dvld[37][OW_DVLD_W-1:0]),
    `endif
        .s37i_data(stream_in_data[37][`STREAM37_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM37_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s37o_rdy(stream_out_rdy[37]),
        .s37o_valid(stream_out_valid[37]),
    `ifdef STREAM37_OUT_256BIT
	.s37o_ow_dvld(stream_out_ow_dvld[37][OW_DVLD_W-1:0]),
    `endif
        .s37o_data(stream_out_data[37][`STREAM37_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM38_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s38i_rdy(stream_in_rdy[38]),
        .s38i_valid(stream_in_valid[38]),
    `ifdef STREAM38_IN_256BIT
	.s38i_ow_dvld(stream_in_ow_dvld[38][OW_DVLD_W-1:0]),
    `endif
        .s38i_data(stream_in_data[38][`STREAM38_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM38_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s38o_rdy(stream_out_rdy[38]),
        .s38o_valid(stream_out_valid[38]),
    `ifdef STREAM38_OUT_256BIT
	.s38o_ow_dvld(stream_out_ow_dvld[38][OW_DVLD_W-1:0]),
    `endif
        .s38o_data(stream_out_data[38][`STREAM38_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM39_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s39i_rdy(stream_in_rdy[39]),
        .s39i_valid(stream_in_valid[39]),
    `ifdef STREAM39_IN_256BIT
	.s39i_ow_dvld(stream_in_ow_dvld[39][OW_DVLD_W-1:0]),
    `endif
        .s39i_data(stream_in_data[39][`STREAM39_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM39_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s39o_rdy(stream_out_rdy[39]),
        .s39o_valid(stream_out_valid[39]),
    `ifdef STREAM39_OUT_256BIT
	.s39o_ow_dvld(stream_out_ow_dvld[39][OW_DVLD_W-1:0]),
    `endif
        .s39o_data(stream_out_data[39][`STREAM39_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM40_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s40i_rdy(stream_in_rdy[40]),
        .s40i_valid(stream_in_valid[40]),
    `ifdef STREAM40_IN_256BIT
	.s40i_ow_dvld(stream_in_ow_dvld[40][OW_DVLD_W-1:0]),
    `endif
        .s40i_data(stream_in_data[40][`STREAM40_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM40_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s40o_rdy(stream_out_rdy[40]),
        .s40o_valid(stream_out_valid[40]),
    `ifdef STREAM40_OUT_256BIT
	.s40o_ow_dvld(stream_out_ow_dvld[40][OW_DVLD_W-1:0]),
    `endif
        .s40o_data(stream_out_data[40][`STREAM40_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM41_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s41i_rdy(stream_in_rdy[41]),
        .s41i_valid(stream_in_valid[41]),
    `ifdef STREAM41_IN_256BIT
	.s41i_ow_dvld(stream_in_ow_dvld[41][OW_DVLD_W-1:0]),
    `endif
        .s41i_data(stream_in_data[41][`STREAM41_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM41_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s41o_rdy(stream_out_rdy[41]),
        .s41o_valid(stream_out_valid[41]),
    `ifdef STREAM41_OUT_256BIT
	.s41o_ow_dvld(stream_out_ow_dvld[41][OW_DVLD_W-1:0]),
    `endif
        .s41o_data(stream_out_data[41][`STREAM41_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM42_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s42i_rdy(stream_in_rdy[42]),
        .s42i_valid(stream_in_valid[42]),
    `ifdef STREAM42_IN_256BIT
	.s42i_ow_dvld(stream_in_ow_dvld[42][OW_DVLD_W-1:0]),
    `endif
        .s42i_data(stream_in_data[42][`STREAM42_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM42_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s42o_rdy(stream_out_rdy[42]),
        .s42o_valid(stream_out_valid[42]),
    `ifdef STREAM42_OUT_256BIT
	.s42o_ow_dvld(stream_out_ow_dvld[42][OW_DVLD_W-1:0]),
    `endif
        .s42o_data(stream_out_data[42][`STREAM42_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM43_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s43i_rdy(stream_in_rdy[43]),
        .s43i_valid(stream_in_valid[43]),
    `ifdef STREAM43_IN_256BIT
	.s43i_ow_dvld(stream_in_ow_dvld[43][OW_DVLD_W-1:0]),
    `endif
        .s43i_data(stream_in_data[43][`STREAM43_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM43_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s43o_rdy(stream_out_rdy[43]),
        .s43o_valid(stream_out_valid[43]),
    `ifdef STREAM43_OUT_256BIT
	.s43o_ow_dvld(stream_out_ow_dvld[43][OW_DVLD_W-1:0]),
    `endif
        .s43o_data(stream_out_data[43][`STREAM43_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM44_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s44i_rdy(stream_in_rdy[44]),
        .s44i_valid(stream_in_valid[44]),
    `ifdef STREAM44_IN_256BIT
	.s44i_ow_dvld(stream_in_ow_dvld[44][OW_DVLD_W-1:0]),
    `endif
        .s44i_data(stream_in_data[44][`STREAM44_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM44_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s44o_rdy(stream_out_rdy[44]),
        .s44o_valid(stream_out_valid[44]),
    `ifdef STREAM44_OUT_256BIT
	.s44o_ow_dvld(stream_out_ow_dvld[44][OW_DVLD_W-1:0]),
    `endif
        .s44o_data(stream_out_data[44][`STREAM44_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM45_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s45i_rdy(stream_in_rdy[45]),
        .s45i_valid(stream_in_valid[45]),
    `ifdef STREAM45_IN_256BIT
	.s45i_ow_dvld(stream_in_ow_dvld[45][OW_DVLD_W-1:0]),
    `endif
        .s45i_data(stream_in_data[45][`STREAM45_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM45_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s45o_rdy(stream_out_rdy[45]),
        .s45o_valid(stream_out_valid[45]),
    `ifdef STREAM45_OUT_256BIT
	.s45o_ow_dvld(stream_out_ow_dvld[45][OW_DVLD_W-1:0]),
    `endif
        .s45o_data(stream_out_data[45][`STREAM45_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM46_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s46i_rdy(stream_in_rdy[46]),
        .s46i_valid(stream_in_valid[46]),
    `ifdef STREAM46_IN_256BIT
	.s46i_ow_dvld(stream_in_ow_dvld[46][OW_DVLD_W-1:0]),
    `endif
        .s46i_data(stream_in_data[46][`STREAM46_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM46_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s46o_rdy(stream_out_rdy[46]),
        .s46o_valid(stream_out_valid[46]),
    `ifdef STREAM46_OUT_256BIT
	.s46o_ow_dvld(stream_out_ow_dvld[46][OW_DVLD_W-1:0]),
    `endif
        .s46o_data(stream_out_data[46][`STREAM46_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM47_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s47i_rdy(stream_in_rdy[47]),
        .s47i_valid(stream_in_valid[47]),
    `ifdef STREAM47_IN_256BIT
	.s47i_ow_dvld(stream_in_ow_dvld[47][OW_DVLD_W-1:0]),
    `endif
        .s47i_data(stream_in_data[47][`STREAM47_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM47_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s47o_rdy(stream_out_rdy[47]),
        .s47o_valid(stream_out_valid[47]),
    `ifdef STREAM47_OUT_256BIT
	.s47o_ow_dvld(stream_out_ow_dvld[47][OW_DVLD_W-1:0]),
    `endif
        .s47o_data(stream_out_data[47][`STREAM47_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM48_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s48i_rdy(stream_in_rdy[48]),
        .s48i_valid(stream_in_valid[48]),
    `ifdef STREAM48_IN_256BIT
	.s48i_ow_dvld(stream_in_ow_dvld[48][OW_DVLD_W-1:0]),
    `endif
        .s48i_data(stream_in_data[48][`STREAM48_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM48_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s48o_rdy(stream_out_rdy[48]),
        .s48o_valid(stream_out_valid[48]),
    `ifdef STREAM48_OUT_256BIT
	.s48o_ow_dvld(stream_out_ow_dvld[48][OW_DVLD_W-1:0]),
    `endif
        .s48o_data(stream_out_data[48][`STREAM48_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM49_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s49i_rdy(stream_in_rdy[49]),
        .s49i_valid(stream_in_valid[49]),
    `ifdef STREAM49_IN_256BIT
	.s49i_ow_dvld(stream_in_ow_dvld[49][OW_DVLD_W-1:0]),
    `endif
        .s49i_data(stream_in_data[49][`STREAM49_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM49_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s49o_rdy(stream_out_rdy[49]),
        .s49o_valid(stream_out_valid[49]),
    `ifdef STREAM49_OUT_256BIT
	.s49o_ow_dvld(stream_out_ow_dvld[49][OW_DVLD_W-1:0]),
    `endif
        .s49o_data(stream_out_data[49][`STREAM49_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM50_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s50i_rdy(stream_in_rdy[50]),
        .s50i_valid(stream_in_valid[50]),
    `ifdef STREAM50_IN_256BIT
	.s50i_ow_dvld(stream_in_ow_dvld[50][OW_DVLD_W-1:0]),
    `endif
        .s50i_data(stream_in_data[50][`STREAM50_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM50_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s50o_rdy(stream_out_rdy[50]),
        .s50o_valid(stream_out_valid[50]),
    `ifdef STREAM50_OUT_256BIT
	.s50o_ow_dvld(stream_out_ow_dvld[50][OW_DVLD_W-1:0]),
    `endif
        .s50o_data(stream_out_data[50][`STREAM50_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM51_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s51i_rdy(stream_in_rdy[51]),
        .s51i_valid(stream_in_valid[51]),
    `ifdef STREAM51_IN_256BIT
	.s51i_ow_dvld(stream_in_ow_dvld[51][OW_DVLD_W-1:0]),
    `endif
        .s51i_data(stream_in_data[51][`STREAM51_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM51_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s51o_rdy(stream_out_rdy[51]),
        .s51o_valid(stream_out_valid[51]),
    `ifdef STREAM51_OUT_256BIT
	.s51o_ow_dvld(stream_out_ow_dvld[51][OW_DVLD_W-1:0]),
    `endif
        .s51o_data(stream_out_data[51][`STREAM51_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM52_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s52i_rdy(stream_in_rdy[52]),
        .s52i_valid(stream_in_valid[52]),
    `ifdef STREAM52_IN_256BIT
	.s52i_ow_dvld(stream_in_ow_dvld[52][OW_DVLD_W-1:0]),
    `endif
        .s52i_data(stream_in_data[52][`STREAM52_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM52_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s52o_rdy(stream_out_rdy[52]),
        .s52o_valid(stream_out_valid[52]),
    `ifdef STREAM52_OUT_256BIT
	.s52o_ow_dvld(stream_out_ow_dvld[52][OW_DVLD_W-1:0]),
    `endif
        .s52o_data(stream_out_data[52][`STREAM52_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM53_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s53i_rdy(stream_in_rdy[53]),
        .s53i_valid(stream_in_valid[53]),
    `ifdef STREAM53_IN_256BIT
	.s53i_ow_dvld(stream_in_ow_dvld[53][OW_DVLD_W-1:0]),
    `endif
        .s53i_data(stream_in_data[53][`STREAM53_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM53_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s53o_rdy(stream_out_rdy[53]),
        .s53o_valid(stream_out_valid[53]),
    `ifdef STREAM53_OUT_256BIT
	.s53o_ow_dvld(stream_out_ow_dvld[53][OW_DVLD_W-1:0]),
    `endif
        .s53o_data(stream_out_data[53][`STREAM53_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM54_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s54i_rdy(stream_in_rdy[54]),
        .s54i_valid(stream_in_valid[54]),
    `ifdef STREAM54_IN_256BIT
	.s54i_ow_dvld(stream_in_ow_dvld[54][OW_DVLD_W-1:0]),
    `endif
        .s54i_data(stream_in_data[54][`STREAM54_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM54_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s54o_rdy(stream_out_rdy[54]),
        .s54o_valid(stream_out_valid[54]),
    `ifdef STREAM54_OUT_256BIT
	.s54o_ow_dvld(stream_out_ow_dvld[54][OW_DVLD_W-1:0]),
    `endif
        .s54o_data(stream_out_data[54][`STREAM54_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM55_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s55i_rdy(stream_in_rdy[55]),
        .s55i_valid(stream_in_valid[55]),
    `ifdef STREAM55_IN_256BIT
	.s55i_ow_dvld(stream_in_ow_dvld[55][OW_DVLD_W-1:0]),
    `endif
        .s55i_data(stream_in_data[55][`STREAM55_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM55_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s55o_rdy(stream_out_rdy[55]),
        .s55o_valid(stream_out_valid[55]),
    `ifdef STREAM55_OUT_256BIT
	.s55o_ow_dvld(stream_out_ow_dvld[55][OW_DVLD_W-1:0]),
    `endif
        .s55o_data(stream_out_data[55][`STREAM55_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM56_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s56i_rdy(stream_in_rdy[56]),
        .s56i_valid(stream_in_valid[56]),
    `ifdef STREAM56_IN_256BIT
	.s56i_ow_dvld(stream_in_ow_dvld[56][OW_DVLD_W-1:0]),
    `endif
        .s56i_data(stream_in_data[56][`STREAM56_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM56_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s56o_rdy(stream_out_rdy[56]),
        .s56o_valid(stream_out_valid[56]),
    `ifdef STREAM56_OUT_256BIT
	.s56o_ow_dvld(stream_out_ow_dvld[56][OW_DVLD_W-1:0]),
    `endif
        .s56o_data(stream_out_data[56][`STREAM56_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM57_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s57i_rdy(stream_in_rdy[57]),
        .s57i_valid(stream_in_valid[57]),
    `ifdef STREAM57_IN_256BIT
	.s57i_ow_dvld(stream_in_ow_dvld[57][OW_DVLD_W-1:0]),
    `endif
        .s57i_data(stream_in_data[57][`STREAM57_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM57_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s57o_rdy(stream_out_rdy[57]),
        .s57o_valid(stream_out_valid[57]),
    `ifdef STREAM57_OUT_256BIT
	.s57o_ow_dvld(stream_out_ow_dvld[57][OW_DVLD_W-1:0]),
    `endif
        .s57o_data(stream_out_data[57][`STREAM57_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM58_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s58i_rdy(stream_in_rdy[58]),
        .s58i_valid(stream_in_valid[58]),
    `ifdef STREAM58_IN_256BIT
	.s58i_ow_dvld(stream_in_ow_dvld[58][OW_DVLD_W-1:0]),
    `endif
        .s58i_data(stream_in_data[58][`STREAM58_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM58_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s58o_rdy(stream_out_rdy[58]),
        .s58o_valid(stream_out_valid[58]),
    `ifdef STREAM58_OUT_256BIT
	.s58o_ow_dvld(stream_out_ow_dvld[58][OW_DVLD_W-1:0]),
    `endif
        .s58o_data(stream_out_data[58][`STREAM58_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM59_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s59i_rdy(stream_in_rdy[59]),
        .s59i_valid(stream_in_valid[59]),
    `ifdef STREAM59_IN_256BIT
	.s59i_ow_dvld(stream_in_ow_dvld[59][OW_DVLD_W-1:0]),
    `endif
        .s59i_data(stream_in_data[59][`STREAM59_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM59_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s59o_rdy(stream_out_rdy[59]),
        .s59o_valid(stream_out_valid[59]),
    `ifdef STREAM59_OUT_256BIT
	.s59o_ow_dvld(stream_out_ow_dvld[59][OW_DVLD_W-1:0]),
    `endif
        .s59o_data(stream_out_data[59][`STREAM59_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM60_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s60i_rdy(stream_in_rdy[60]),
        .s60i_valid(stream_in_valid[60]),
    `ifdef STREAM60_IN_256BIT
	.s60i_ow_dvld(stream_in_ow_dvld[60][OW_DVLD_W-1:0]),
    `endif
        .s60i_data(stream_in_data[60][`STREAM60_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM60_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s60o_rdy(stream_out_rdy[60]),
        .s60o_valid(stream_out_valid[60]),
    `ifdef STREAM60_OUT_256BIT
	.s60o_ow_dvld(stream_out_ow_dvld[60][OW_DVLD_W-1:0]),
    `endif
        .s60o_data(stream_out_data[60][`STREAM60_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM61_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s61i_rdy(stream_in_rdy[61]),
        .s61i_valid(stream_in_valid[61]),
    `ifdef STREAM61_IN_256BIT
	.s61i_ow_dvld(stream_in_ow_dvld[61][OW_DVLD_W-1:0]),
    `endif
        .s61i_data(stream_in_data[61][`STREAM61_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM61_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s61o_rdy(stream_out_rdy[61]),
        .s61o_valid(stream_out_valid[61]),
    `ifdef STREAM61_OUT_256BIT
	.s61o_ow_dvld(stream_out_ow_dvld[61][OW_DVLD_W-1:0]),
    `endif
        .s61o_data(stream_out_data[61][`STREAM61_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM62_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s62i_rdy(stream_in_rdy[62]),
        .s62i_valid(stream_in_valid[62]),
    `ifdef STREAM62_IN_256BIT
	.s62i_ow_dvld(stream_in_ow_dvld[62][OW_DVLD_W-1:0]),
    `endif
        .s62i_data(stream_in_data[62][`STREAM62_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM62_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s62o_rdy(stream_out_rdy[62]),
        .s62o_valid(stream_out_valid[62]),
    `ifdef STREAM62_OUT_256BIT
	.s62o_ow_dvld(stream_out_ow_dvld[62][OW_DVLD_W-1:0]),
    `endif
        .s62o_data(stream_out_data[62][`STREAM62_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM63_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s63i_rdy(stream_in_rdy[63]),
        .s63i_valid(stream_in_valid[63]),
    `ifdef STREAM63_IN_256BIT
	.s63i_ow_dvld(stream_in_ow_dvld[63][OW_DVLD_W-1:0]),
    `endif
        .s63i_data(stream_in_data[63][`STREAM63_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM63_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s63o_rdy(stream_out_rdy[63]),
        .s63o_valid(stream_out_valid[63]),
    `ifdef STREAM63_OUT_256BIT
	.s63o_ow_dvld(stream_out_ow_dvld[63][OW_DVLD_W-1:0]),
    `endif
        .s63o_data(stream_out_data[63][`STREAM63_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM64_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s64i_rdy(stream_in_rdy[64]),
        .s64i_valid(stream_in_valid[64]),
    `ifdef STREAM64_IN_256BIT
	.s64i_ow_dvld(stream_in_ow_dvld[64][OW_DVLD_W-1:0]),
    `endif
        .s64i_data(stream_in_data[64][`STREAM64_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM64_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s64o_rdy(stream_out_rdy[64]),
        .s64o_valid(stream_out_valid[64]),
    `ifdef STREAM64_OUT_256BIT
	.s64o_ow_dvld(stream_out_ow_dvld[64][OW_DVLD_W-1:0]),
    `endif
        .s64o_data(stream_out_data[64][`STREAM64_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM65_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s65i_rdy(stream_in_rdy[65]),
        .s65i_valid(stream_in_valid[65]),
    `ifdef STREAM65_IN_256BIT
	.s65i_ow_dvld(stream_in_ow_dvld[65][OW_DVLD_W-1:0]),
    `endif
        .s65i_data(stream_in_data[65][`STREAM65_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM65_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s65o_rdy(stream_out_rdy[65]),
        .s65o_valid(stream_out_valid[65]),
    `ifdef STREAM65_OUT_256BIT
	.s65o_ow_dvld(stream_out_ow_dvld[65][OW_DVLD_W-1:0]),
    `endif
        .s65o_data(stream_out_data[65][`STREAM65_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM66_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s66i_rdy(stream_in_rdy[66]),
        .s66i_valid(stream_in_valid[66]),
    `ifdef STREAM66_IN_256BIT
	.s66i_ow_dvld(stream_in_ow_dvld[66][OW_DVLD_W-1:0]),
    `endif
        .s66i_data(stream_in_data[66][`STREAM66_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM66_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s66o_rdy(stream_out_rdy[66]),
        .s66o_valid(stream_out_valid[66]),
    `ifdef STREAM66_OUT_256BIT
	.s66o_ow_dvld(stream_out_ow_dvld[66][OW_DVLD_W-1:0]),
    `endif
        .s66o_data(stream_out_data[66][`STREAM66_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM67_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s67i_rdy(stream_in_rdy[67]),
        .s67i_valid(stream_in_valid[67]),
    `ifdef STREAM67_IN_256BIT
	.s67i_ow_dvld(stream_in_ow_dvld[67][OW_DVLD_W-1:0]),
    `endif
        .s67i_data(stream_in_data[67][`STREAM67_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM67_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s67o_rdy(stream_out_rdy[67]),
        .s67o_valid(stream_out_valid[67]),
    `ifdef STREAM67_OUT_256BIT
	.s67o_ow_dvld(stream_out_ow_dvld[67][OW_DVLD_W-1:0]),
    `endif
        .s67o_data(stream_out_data[67][`STREAM67_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM68_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s68i_rdy(stream_in_rdy[68]),
        .s68i_valid(stream_in_valid[68]),
    `ifdef STREAM68_IN_256BIT
	.s68i_ow_dvld(stream_in_ow_dvld[68][OW_DVLD_W-1:0]),
    `endif
        .s68i_data(stream_in_data[68][`STREAM68_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM68_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s68o_rdy(stream_out_rdy[68]),
        .s68o_valid(stream_out_valid[68]),
    `ifdef STREAM68_OUT_256BIT
	.s68o_ow_dvld(stream_out_ow_dvld[68][OW_DVLD_W-1:0]),
    `endif
        .s68o_data(stream_out_data[68][`STREAM68_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM69_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s69i_rdy(stream_in_rdy[69]),
        .s69i_valid(stream_in_valid[69]),
    `ifdef STREAM69_IN_256BIT
	.s69i_ow_dvld(stream_in_ow_dvld[69][OW_DVLD_W-1:0]),
    `endif
        .s69i_data(stream_in_data[69][`STREAM69_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM69_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s69o_rdy(stream_out_rdy[69]),
        .s69o_valid(stream_out_valid[69]),
    `ifdef STREAM69_OUT_256BIT
	.s69o_ow_dvld(stream_out_ow_dvld[69][OW_DVLD_W-1:0]),
    `endif
        .s69o_data(stream_out_data[69][`STREAM69_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM70_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s70i_rdy(stream_in_rdy[70]),
        .s70i_valid(stream_in_valid[70]),
    `ifdef STREAM70_IN_256BIT
	.s70i_ow_dvld(stream_in_ow_dvld[70][OW_DVLD_W-1:0]),
    `endif
        .s70i_data(stream_in_data[70][`STREAM70_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM70_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s70o_rdy(stream_out_rdy[70]),
        .s70o_valid(stream_out_valid[70]),
    `ifdef STREAM70_OUT_256BIT
	.s70o_ow_dvld(stream_out_ow_dvld[70][OW_DVLD_W-1:0]),
    `endif
        .s70o_data(stream_out_data[70][`STREAM70_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM71_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s71i_rdy(stream_in_rdy[71]),
        .s71i_valid(stream_in_valid[71]),
    `ifdef STREAM71_IN_256BIT
	.s71i_ow_dvld(stream_in_ow_dvld[71][OW_DVLD_W-1:0]),
    `endif
        .s71i_data(stream_in_data[71][`STREAM71_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM71_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s71o_rdy(stream_out_rdy[71]),
        .s71o_valid(stream_out_valid[71]),
    `ifdef STREAM71_OUT_256BIT
	.s71o_ow_dvld(stream_out_ow_dvld[71][OW_DVLD_W-1:0]),
    `endif
        .s71o_data(stream_out_data[71][`STREAM71_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM72_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s72i_rdy(stream_in_rdy[72]),
        .s72i_valid(stream_in_valid[72]),
    `ifdef STREAM72_IN_256BIT
	.s72i_ow_dvld(stream_in_ow_dvld[72][OW_DVLD_W-1:0]),
    `endif
        .s72i_data(stream_in_data[72][`STREAM72_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM72_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s72o_rdy(stream_out_rdy[72]),
        .s72o_valid(stream_out_valid[72]),
    `ifdef STREAM72_OUT_256BIT
	.s72o_ow_dvld(stream_out_ow_dvld[72][OW_DVLD_W-1:0]),
    `endif
        .s72o_data(stream_out_data[72][`STREAM72_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM73_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s73i_rdy(stream_in_rdy[73]),
        .s73i_valid(stream_in_valid[73]),
    `ifdef STREAM73_IN_256BIT
	.s73i_ow_dvld(stream_in_ow_dvld[73][OW_DVLD_W-1:0]),
    `endif
        .s73i_data(stream_in_data[73][`STREAM73_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM73_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s73o_rdy(stream_out_rdy[73]),
        .s73o_valid(stream_out_valid[73]),
    `ifdef STREAM73_OUT_256BIT
	.s73o_ow_dvld(stream_out_ow_dvld[73][OW_DVLD_W-1:0]),
    `endif
        .s73o_data(stream_out_data[73][`STREAM73_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM74_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s74i_rdy(stream_in_rdy[74]),
        .s74i_valid(stream_in_valid[74]),
    `ifdef STREAM74_IN_256BIT
	.s74i_ow_dvld(stream_in_ow_dvld[74][OW_DVLD_W-1:0]),
    `endif
        .s74i_data(stream_in_data[74][`STREAM74_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM74_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s74o_rdy(stream_out_rdy[74]),
        .s74o_valid(stream_out_valid[74]),
    `ifdef STREAM74_OUT_256BIT
	.s74o_ow_dvld(stream_out_ow_dvld[74][OW_DVLD_W-1:0]),
    `endif
        .s74o_data(stream_out_data[74][`STREAM74_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM75_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s75i_rdy(stream_in_rdy[75]),
        .s75i_valid(stream_in_valid[75]),
    `ifdef STREAM75_IN_256BIT
	.s75i_ow_dvld(stream_in_ow_dvld[75][OW_DVLD_W-1:0]),
    `endif
        .s75i_data(stream_in_data[75][`STREAM75_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM75_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s75o_rdy(stream_out_rdy[75]),
        .s75o_valid(stream_out_valid[75]),
    `ifdef STREAM75_OUT_256BIT
	.s75o_ow_dvld(stream_out_ow_dvld[75][OW_DVLD_W-1:0]),
    `endif
        .s75o_data(stream_out_data[75][`STREAM75_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM76_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s76i_rdy(stream_in_rdy[76]),
        .s76i_valid(stream_in_valid[76]),
    `ifdef STREAM76_IN_256BIT
	.s76i_ow_dvld(stream_in_ow_dvld[76][OW_DVLD_W-1:0]),
    `endif
        .s76i_data(stream_in_data[76][`STREAM76_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM76_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s76o_rdy(stream_out_rdy[76]),
        .s76o_valid(stream_out_valid[76]),
    `ifdef STREAM76_OUT_256BIT
	.s76o_ow_dvld(stream_out_ow_dvld[76][OW_DVLD_W-1:0]),
    `endif
        .s76o_data(stream_out_data[76][`STREAM76_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM77_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s77i_rdy(stream_in_rdy[77]),
        .s77i_valid(stream_in_valid[77]),
    `ifdef STREAM77_IN_256BIT
	.s77i_ow_dvld(stream_in_ow_dvld[77][OW_DVLD_W-1:0]),
    `endif
        .s77i_data(stream_in_data[77][`STREAM77_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM77_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s77o_rdy(stream_out_rdy[77]),
        .s77o_valid(stream_out_valid[77]),
    `ifdef STREAM77_OUT_256BIT
	.s77o_ow_dvld(stream_out_ow_dvld[77][OW_DVLD_W-1:0]),
    `endif
        .s77o_data(stream_out_data[77][`STREAM77_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM78_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s78i_rdy(stream_in_rdy[78]),
        .s78i_valid(stream_in_valid[78]),
    `ifdef STREAM78_IN_256BIT
	.s78i_ow_dvld(stream_in_ow_dvld[78][OW_DVLD_W-1:0]),
    `endif
        .s78i_data(stream_in_data[78][`STREAM78_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM78_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s78o_rdy(stream_out_rdy[78]),
        .s78o_valid(stream_out_valid[78]),
    `ifdef STREAM78_OUT_256BIT
	.s78o_ow_dvld(stream_out_ow_dvld[78][OW_DVLD_W-1:0]),
    `endif
        .s78o_data(stream_out_data[78][`STREAM78_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM79_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s79i_rdy(stream_in_rdy[79]),
        .s79i_valid(stream_in_valid[79]),
    `ifdef STREAM79_IN_256BIT
	.s79i_ow_dvld(stream_in_ow_dvld[79][OW_DVLD_W-1:0]),
    `endif
        .s79i_data(stream_in_data[79][`STREAM79_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM79_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s79o_rdy(stream_out_rdy[79]),
        .s79o_valid(stream_out_valid[79]),
    `ifdef STREAM79_OUT_256BIT
	.s79o_ow_dvld(stream_out_ow_dvld[79][OW_DVLD_W-1:0]),
    `endif
        .s79o_data(stream_out_data[79][`STREAM79_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM80_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s80i_rdy(stream_in_rdy[80]),
        .s80i_valid(stream_in_valid[80]),
    `ifdef STREAM80_IN_256BIT
	.s80i_ow_dvld(stream_in_ow_dvld[80][OW_DVLD_W-1:0]),
    `endif
        .s80i_data(stream_in_data[80][`STREAM80_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM80_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s80o_rdy(stream_out_rdy[80]),
        .s80o_valid(stream_out_valid[80]),
    `ifdef STREAM80_OUT_256BIT
	.s80o_ow_dvld(stream_out_ow_dvld[80][OW_DVLD_W-1:0]),
    `endif
        .s80o_data(stream_out_data[80][`STREAM80_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM81_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s81i_rdy(stream_in_rdy[81]),
        .s81i_valid(stream_in_valid[81]),
    `ifdef STREAM81_IN_256BIT
	.s81i_ow_dvld(stream_in_ow_dvld[81][OW_DVLD_W-1:0]),
    `endif
        .s81i_data(stream_in_data[81][`STREAM81_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM81_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s81o_rdy(stream_out_rdy[81]),
        .s81o_valid(stream_out_valid[81]),
    `ifdef STREAM81_OUT_256BIT
	.s81o_ow_dvld(stream_out_ow_dvld[81][OW_DVLD_W-1:0]),
    `endif
        .s81o_data(stream_out_data[81][`STREAM81_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM82_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s82i_rdy(stream_in_rdy[82]),
        .s82i_valid(stream_in_valid[82]),
    `ifdef STREAM82_IN_256BIT
	.s82i_ow_dvld(stream_in_ow_dvld[82][OW_DVLD_W-1:0]),
    `endif
        .s82i_data(stream_in_data[82][`STREAM82_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM82_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s82o_rdy(stream_out_rdy[82]),
        .s82o_valid(stream_out_valid[82]),
    `ifdef STREAM82_OUT_256BIT
	.s82o_ow_dvld(stream_out_ow_dvld[82][OW_DVLD_W-1:0]),
    `endif
        .s82o_data(stream_out_data[82][`STREAM82_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM83_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s83i_rdy(stream_in_rdy[83]),
        .s83i_valid(stream_in_valid[83]),
    `ifdef STREAM83_IN_256BIT
	.s83i_ow_dvld(stream_in_ow_dvld[83][OW_DVLD_W-1:0]),
    `endif
        .s83i_data(stream_in_data[83][`STREAM83_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM83_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s83o_rdy(stream_out_rdy[83]),
        .s83o_valid(stream_out_valid[83]),
    `ifdef STREAM83_OUT_256BIT
	.s83o_ow_dvld(stream_out_ow_dvld[83][OW_DVLD_W-1:0]),
    `endif
        .s83o_data(stream_out_data[83][`STREAM83_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM84_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s84i_rdy(stream_in_rdy[84]),
        .s84i_valid(stream_in_valid[84]),
    `ifdef STREAM84_IN_256BIT
	.s84i_ow_dvld(stream_in_ow_dvld[84][OW_DVLD_W-1:0]),
    `endif
        .s84i_data(stream_in_data[84][`STREAM84_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM84_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s84o_rdy(stream_out_rdy[84]),
        .s84o_valid(stream_out_valid[84]),
    `ifdef STREAM84_OUT_256BIT
	.s84o_ow_dvld(stream_out_ow_dvld[84][OW_DVLD_W-1:0]),
    `endif
        .s84o_data(stream_out_data[84][`STREAM84_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM85_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s85i_rdy(stream_in_rdy[85]),
        .s85i_valid(stream_in_valid[85]),
    `ifdef STREAM85_IN_256BIT
	.s85i_ow_dvld(stream_in_ow_dvld[85][OW_DVLD_W-1:0]),
    `endif
        .s85i_data(stream_in_data[85][`STREAM85_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM85_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s85o_rdy(stream_out_rdy[85]),
        .s85o_valid(stream_out_valid[85]),
    `ifdef STREAM85_OUT_256BIT
	.s85o_ow_dvld(stream_out_ow_dvld[85][OW_DVLD_W-1:0]),
    `endif
        .s85o_data(stream_out_data[85][`STREAM85_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM86_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s86i_rdy(stream_in_rdy[86]),
        .s86i_valid(stream_in_valid[86]),
    `ifdef STREAM86_IN_256BIT
	.s86i_ow_dvld(stream_in_ow_dvld[86][OW_DVLD_W-1:0]),
    `endif
        .s86i_data(stream_in_data[86][`STREAM86_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM86_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s86o_rdy(stream_out_rdy[86]),
        .s86o_valid(stream_out_valid[86]),
    `ifdef STREAM86_OUT_256BIT
	.s86o_ow_dvld(stream_out_ow_dvld[86][OW_DVLD_W-1:0]),
    `endif
        .s86o_data(stream_out_data[86][`STREAM86_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM87_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s87i_rdy(stream_in_rdy[87]),
        .s87i_valid(stream_in_valid[87]),
    `ifdef STREAM87_IN_256BIT
	.s87i_ow_dvld(stream_in_ow_dvld[87][OW_DVLD_W-1:0]),
    `endif
        .s87i_data(stream_in_data[87][`STREAM87_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM87_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s87o_rdy(stream_out_rdy[87]),
        .s87o_valid(stream_out_valid[87]),
    `ifdef STREAM87_OUT_256BIT
	.s87o_ow_dvld(stream_out_ow_dvld[87][OW_DVLD_W-1:0]),
    `endif
        .s87o_data(stream_out_data[87][`STREAM87_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM88_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s88i_rdy(stream_in_rdy[88]),
        .s88i_valid(stream_in_valid[88]),
    `ifdef STREAM88_IN_256BIT
	.s88i_ow_dvld(stream_in_ow_dvld[88][OW_DVLD_W-1:0]),
    `endif
        .s88i_data(stream_in_data[88][`STREAM88_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM88_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s88o_rdy(stream_out_rdy[88]),
        .s88o_valid(stream_out_valid[88]),
    `ifdef STREAM88_OUT_256BIT
	.s88o_ow_dvld(stream_out_ow_dvld[88][OW_DVLD_W-1:0]),
    `endif
        .s88o_data(stream_out_data[88][`STREAM88_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM89_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s89i_rdy(stream_in_rdy[89]),
        .s89i_valid(stream_in_valid[89]),
    `ifdef STREAM89_IN_256BIT
	.s89i_ow_dvld(stream_in_ow_dvld[89][OW_DVLD_W-1:0]),
    `endif
        .s89i_data(stream_in_data[89][`STREAM89_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM89_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s89o_rdy(stream_out_rdy[89]),
        .s89o_valid(stream_out_valid[89]),
    `ifdef STREAM89_OUT_256BIT
	.s89o_ow_dvld(stream_out_ow_dvld[89][OW_DVLD_W-1:0]),
    `endif
        .s89o_data(stream_out_data[89][`STREAM89_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM90_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s90i_rdy(stream_in_rdy[90]),
        .s90i_valid(stream_in_valid[90]),
    `ifdef STREAM90_IN_256BIT
	.s90i_ow_dvld(stream_in_ow_dvld[90][OW_DVLD_W-1:0]),
    `endif
        .s90i_data(stream_in_data[90][`STREAM90_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM90_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s90o_rdy(stream_out_rdy[90]),
        .s90o_valid(stream_out_valid[90]),
    `ifdef STREAM90_OUT_256BIT
	.s90o_ow_dvld(stream_out_ow_dvld[90][OW_DVLD_W-1:0]),
    `endif
        .s90o_data(stream_out_data[90][`STREAM90_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM91_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s91i_rdy(stream_in_rdy[91]),
        .s91i_valid(stream_in_valid[91]),
    `ifdef STREAM91_IN_256BIT
	.s91i_ow_dvld(stream_in_ow_dvld[91][OW_DVLD_W-1:0]),
    `endif
        .s91i_data(stream_in_data[91][`STREAM91_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM91_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s91o_rdy(stream_out_rdy[91]),
        .s91o_valid(stream_out_valid[91]),
    `ifdef STREAM91_OUT_256BIT
	.s91o_ow_dvld(stream_out_ow_dvld[91][OW_DVLD_W-1:0]),
    `endif
        .s91o_data(stream_out_data[91][`STREAM91_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM92_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s92i_rdy(stream_in_rdy[92]),
        .s92i_valid(stream_in_valid[92]),
    `ifdef STREAM92_IN_256BIT
	.s92i_ow_dvld(stream_in_ow_dvld[92][OW_DVLD_W-1:0]),
    `endif
        .s92i_data(stream_in_data[92][`STREAM92_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM92_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s92o_rdy(stream_out_rdy[92]),
        .s92o_valid(stream_out_valid[92]),
    `ifdef STREAM92_OUT_256BIT
	.s92o_ow_dvld(stream_out_ow_dvld[92][OW_DVLD_W-1:0]),
    `endif
        .s92o_data(stream_out_data[92][`STREAM92_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM93_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s93i_rdy(stream_in_rdy[93]),
        .s93i_valid(stream_in_valid[93]),
    `ifdef STREAM93_IN_256BIT
	.s93i_ow_dvld(stream_in_ow_dvld[93][OW_DVLD_W-1:0]),
    `endif
        .s93i_data(stream_in_data[93][`STREAM93_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM93_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s93o_rdy(stream_out_rdy[93]),
        .s93o_valid(stream_out_valid[93]),
    `ifdef STREAM93_OUT_256BIT
	.s93o_ow_dvld(stream_out_ow_dvld[93][OW_DVLD_W-1:0]),
    `endif
        .s93o_data(stream_out_data[93][`STREAM93_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM94_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s94i_rdy(stream_in_rdy[94]),
        .s94i_valid(stream_in_valid[94]),
    `ifdef STREAM94_IN_256BIT
	.s94i_ow_dvld(stream_in_ow_dvld[94][OW_DVLD_W-1:0]),
    `endif
        .s94i_data(stream_in_data[94][`STREAM94_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM94_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s94o_rdy(stream_out_rdy[94]),
        .s94o_valid(stream_out_valid[94]),
    `ifdef STREAM94_OUT_256BIT
	.s94o_ow_dvld(stream_out_ow_dvld[94][OW_DVLD_W-1:0]),
    `endif
        .s94o_data(stream_out_data[94][`STREAM94_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM95_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s95i_rdy(stream_in_rdy[95]),
        .s95i_valid(stream_in_valid[95]),
    `ifdef STREAM95_IN_256BIT
	.s95i_ow_dvld(stream_in_ow_dvld[95][OW_DVLD_W-1:0]),
    `endif
        .s95i_data(stream_in_data[95][`STREAM95_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM95_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s95o_rdy(stream_out_rdy[95]),
        .s95o_valid(stream_out_valid[95]),
    `ifdef STREAM95_OUT_256BIT
	.s95o_ow_dvld(stream_out_ow_dvld[95][OW_DVLD_W-1:0]),
    `endif
        .s95o_data(stream_out_data[95][`STREAM95_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM96_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s96i_rdy(stream_in_rdy[96]),
        .s96i_valid(stream_in_valid[96]),
    `ifdef STREAM96_IN_256BIT
	.s96i_ow_dvld(stream_in_ow_dvld[96][OW_DVLD_W-1:0]),
    `endif
        .s96i_data(stream_in_data[96][`STREAM96_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM96_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s96o_rdy(stream_out_rdy[96]),
        .s96o_valid(stream_out_valid[96]),
    `ifdef STREAM96_OUT_256BIT
	.s96o_ow_dvld(stream_out_ow_dvld[96][OW_DVLD_W-1:0]),
    `endif
        .s96o_data(stream_out_data[96][`STREAM96_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM97_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s97i_rdy(stream_in_rdy[97]),
        .s97i_valid(stream_in_valid[97]),
    `ifdef STREAM97_IN_256BIT
	.s97i_ow_dvld(stream_in_ow_dvld[97][OW_DVLD_W-1:0]),
    `endif
        .s97i_data(stream_in_data[97][`STREAM97_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM97_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s97o_rdy(stream_out_rdy[97]),
        .s97o_valid(stream_out_valid[97]),
    `ifdef STREAM97_OUT_256BIT
	.s97o_ow_dvld(stream_out_ow_dvld[97][OW_DVLD_W-1:0]),
    `endif
        .s97o_data(stream_out_data[97][`STREAM97_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM98_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s98i_rdy(stream_in_rdy[98]),
        .s98i_valid(stream_in_valid[98]),
    `ifdef STREAM98_IN_256BIT
	.s98i_ow_dvld(stream_in_ow_dvld[98][OW_DVLD_W-1:0]),
    `endif
        .s98i_data(stream_in_data[98][`STREAM98_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM98_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s98o_rdy(stream_out_rdy[98]),
        .s98o_valid(stream_out_valid[98]),
    `ifdef STREAM98_OUT_256BIT
	.s98o_ow_dvld(stream_out_ow_dvld[98][OW_DVLD_W-1:0]),
    `endif
        .s98o_data(stream_out_data[98][`STREAM98_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM99_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s99i_rdy(stream_in_rdy[99]),
        .s99i_valid(stream_in_valid[99]),
    `ifdef STREAM99_IN_256BIT
	.s99i_ow_dvld(stream_in_ow_dvld[99][OW_DVLD_W-1:0]),
    `endif
        .s99i_data(stream_in_data[99][`STREAM99_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM99_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s99o_rdy(stream_out_rdy[99]),
        .s99o_valid(stream_out_valid[99]),
    `ifdef STREAM99_OUT_256BIT
	.s99o_ow_dvld(stream_out_ow_dvld[99][OW_DVLD_W-1:0]),
    `endif
        .s99o_data(stream_out_data[99][`STREAM99_OUT_WIDTH-1:0])
    `endif
    `ifdef STREAM100_IN_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s100i_rdy(stream_in_rdy[100]),
        .s100i_valid(stream_in_valid[100]),
    `ifdef STREAM100_IN_256BIT
	.s100i_ow_dvld(stream_in_ow_dvld[100][OW_DVLD_W-1:0]),
    `endif
        .s100i_data(stream_in_data[100][`STREAM100_IN_WIDTH-1:0])
    `endif
    `ifdef STREAM100_OUT_WIDTH
        `ifdef  UM_PREPEND_COMMA , `endif
        `define UM_PREPEND_COMMA
        `define INCLUDE_STREAM_COMMON
        .s100o_rdy(stream_out_rdy[100]),
        .s100o_valid(stream_out_valid[100]),
    `ifdef STREAM100_OUT_256BIT
	.s100o_ow_dvld(stream_out_ow_dvld[100][OW_DVLD_W-1:0]),
    `endif
        .s100o_data(stream_out_data[100][`STREAM100_OUT_WIDTH-1:0])
    `endif
    `undef UM_PREPEND_COMMA

    `ifdef INCLUDE_STREAM_COMMON
        ,.clk(clk),
        .rst(rst)
    `endif

    );
`endif

// This is the stream compression for the in and out streams into the single signal which is transmited back across to the host.

    assign s_poll_seq[31:0]         = (32'h0
                                        `ifdef PICOBUS_WIDTH  | s_poll_seq_userpb     `endif
                                        `ifdef STREAM1_IN_WIDTH  | stream_in_desc_poll_seq[1]  `endif
                                        `ifdef STREAM1_OUT_WIDTH | stream_out_desc_poll_seq[1] `endif
                                        `ifdef STREAM2_IN_WIDTH  | stream_in_desc_poll_seq[2]  `endif
                                        `ifdef STREAM2_OUT_WIDTH | stream_out_desc_poll_seq[2] `endif
                                        `ifdef STREAM3_IN_WIDTH  | stream_in_desc_poll_seq[3]  `endif
                                        `ifdef STREAM3_OUT_WIDTH | stream_out_desc_poll_seq[3] `endif
                                        `ifdef STREAM4_IN_WIDTH  | stream_in_desc_poll_seq[4]  `endif
                                        `ifdef STREAM4_OUT_WIDTH | stream_out_desc_poll_seq[4] `endif
                                        `ifdef STREAM5_IN_WIDTH  | stream_in_desc_poll_seq[5]  `endif
                                        `ifdef STREAM5_OUT_WIDTH | stream_out_desc_poll_seq[5] `endif
                                        `ifdef STREAM6_IN_WIDTH  | stream_in_desc_poll_seq[6]  `endif
                                        `ifdef STREAM6_OUT_WIDTH | stream_out_desc_poll_seq[6] `endif
                                        `ifdef STREAM7_IN_WIDTH  | stream_in_desc_poll_seq[7]  `endif
                                        `ifdef STREAM7_OUT_WIDTH | stream_out_desc_poll_seq[7] `endif
                                        `ifdef STREAM8_IN_WIDTH  | stream_in_desc_poll_seq[8]  `endif
                                        `ifdef STREAM8_OUT_WIDTH | stream_out_desc_poll_seq[8] `endif
                                        `ifdef STREAM9_IN_WIDTH  | stream_in_desc_poll_seq[9]  `endif
                                        `ifdef STREAM9_OUT_WIDTH | stream_out_desc_poll_seq[9] `endif
                                        `ifdef STREAM10_IN_WIDTH  | stream_in_desc_poll_seq[10]  `endif
                                        `ifdef STREAM10_OUT_WIDTH | stream_out_desc_poll_seq[10] `endif
                                        `ifdef STREAM11_IN_WIDTH  | stream_in_desc_poll_seq[11]  `endif
                                        `ifdef STREAM11_OUT_WIDTH | stream_out_desc_poll_seq[11] `endif
                                        `ifdef STREAM12_IN_WIDTH  | stream_in_desc_poll_seq[12]  `endif
                                        `ifdef STREAM12_OUT_WIDTH | stream_out_desc_poll_seq[12] `endif
                                        `ifdef STREAM13_IN_WIDTH  | stream_in_desc_poll_seq[13]  `endif
                                        `ifdef STREAM13_OUT_WIDTH | stream_out_desc_poll_seq[13] `endif
                                        `ifdef STREAM14_IN_WIDTH  | stream_in_desc_poll_seq[14]  `endif
                                        `ifdef STREAM14_OUT_WIDTH | stream_out_desc_poll_seq[14] `endif
                                        `ifdef STREAM15_IN_WIDTH  | stream_in_desc_poll_seq[15]  `endif
                                        `ifdef STREAM15_OUT_WIDTH | stream_out_desc_poll_seq[15] `endif
                                        `ifdef STREAM16_IN_WIDTH  | stream_in_desc_poll_seq[16]  `endif
                                        `ifdef STREAM16_OUT_WIDTH | stream_out_desc_poll_seq[16] `endif
                                        `ifdef STREAM17_IN_WIDTH  | stream_in_desc_poll_seq[17]  `endif
                                        `ifdef STREAM17_OUT_WIDTH | stream_out_desc_poll_seq[17] `endif
                                        `ifdef STREAM18_IN_WIDTH  | stream_in_desc_poll_seq[18]  `endif
                                        `ifdef STREAM18_OUT_WIDTH | stream_out_desc_poll_seq[18] `endif
                                        `ifdef STREAM19_IN_WIDTH  | stream_in_desc_poll_seq[19]  `endif
                                        `ifdef STREAM19_OUT_WIDTH | stream_out_desc_poll_seq[19] `endif
                                        `ifdef STREAM20_IN_WIDTH  | stream_in_desc_poll_seq[20]  `endif
                                        `ifdef STREAM20_OUT_WIDTH | stream_out_desc_poll_seq[20] `endif
                                        `ifdef STREAM21_IN_WIDTH  | stream_in_desc_poll_seq[21]  `endif
                                        `ifdef STREAM21_OUT_WIDTH | stream_out_desc_poll_seq[21] `endif
                                        `ifdef STREAM22_IN_WIDTH  | stream_in_desc_poll_seq[22]  `endif
                                        `ifdef STREAM22_OUT_WIDTH | stream_out_desc_poll_seq[22] `endif
                                        `ifdef STREAM23_IN_WIDTH  | stream_in_desc_poll_seq[23]  `endif
                                        `ifdef STREAM23_OUT_WIDTH | stream_out_desc_poll_seq[23] `endif
                                        `ifdef STREAM24_IN_WIDTH  | stream_in_desc_poll_seq[24]  `endif
                                        `ifdef STREAM24_OUT_WIDTH | stream_out_desc_poll_seq[24] `endif
                                        `ifdef STREAM25_IN_WIDTH  | stream_in_desc_poll_seq[25]  `endif
                                        `ifdef STREAM25_OUT_WIDTH | stream_out_desc_poll_seq[25] `endif
                                        `ifdef STREAM26_IN_WIDTH  | stream_in_desc_poll_seq[26]  `endif
                                        `ifdef STREAM26_OUT_WIDTH | stream_out_desc_poll_seq[26] `endif
                                        `ifdef STREAM27_IN_WIDTH  | stream_in_desc_poll_seq[27]  `endif
                                        `ifdef STREAM27_OUT_WIDTH | stream_out_desc_poll_seq[27] `endif
                                        `ifdef STREAM28_IN_WIDTH  | stream_in_desc_poll_seq[28]  `endif
                                        `ifdef STREAM28_OUT_WIDTH | stream_out_desc_poll_seq[28] `endif
                                        `ifdef STREAM29_IN_WIDTH  | stream_in_desc_poll_seq[29]  `endif
                                        `ifdef STREAM29_OUT_WIDTH | stream_out_desc_poll_seq[29] `endif
                                        `ifdef STREAM30_IN_WIDTH  | stream_in_desc_poll_seq[30]  `endif
                                        `ifdef STREAM30_OUT_WIDTH | stream_out_desc_poll_seq[30] `endif
                                        `ifdef STREAM31_IN_WIDTH  | stream_in_desc_poll_seq[31]  `endif
                                        `ifdef STREAM31_OUT_WIDTH | stream_out_desc_poll_seq[31] `endif
                                        `ifdef STREAM32_IN_WIDTH  | stream_in_desc_poll_seq[32]  `endif
                                        `ifdef STREAM32_OUT_WIDTH | stream_out_desc_poll_seq[32] `endif
                                        `ifdef STREAM33_IN_WIDTH  | stream_in_desc_poll_seq[33]  `endif
                                        `ifdef STREAM33_OUT_WIDTH | stream_out_desc_poll_seq[33] `endif
                                        `ifdef STREAM34_IN_WIDTH  | stream_in_desc_poll_seq[34]  `endif
                                        `ifdef STREAM34_OUT_WIDTH | stream_out_desc_poll_seq[34] `endif
                                        `ifdef STREAM35_IN_WIDTH  | stream_in_desc_poll_seq[35]  `endif
                                        `ifdef STREAM35_OUT_WIDTH | stream_out_desc_poll_seq[35] `endif
                                        `ifdef STREAM36_IN_WIDTH  | stream_in_desc_poll_seq[36]  `endif
                                        `ifdef STREAM36_OUT_WIDTH | stream_out_desc_poll_seq[36] `endif
                                        `ifdef STREAM37_IN_WIDTH  | stream_in_desc_poll_seq[37]  `endif
                                        `ifdef STREAM37_OUT_WIDTH | stream_out_desc_poll_seq[37] `endif
                                        `ifdef STREAM38_IN_WIDTH  | stream_in_desc_poll_seq[38]  `endif
                                        `ifdef STREAM38_OUT_WIDTH | stream_out_desc_poll_seq[38] `endif
                                        `ifdef STREAM39_IN_WIDTH  | stream_in_desc_poll_seq[39]  `endif
                                        `ifdef STREAM39_OUT_WIDTH | stream_out_desc_poll_seq[39] `endif
                                        `ifdef STREAM40_IN_WIDTH  | stream_in_desc_poll_seq[40]  `endif
                                        `ifdef STREAM40_OUT_WIDTH | stream_out_desc_poll_seq[40] `endif
                                        `ifdef STREAM41_IN_WIDTH  | stream_in_desc_poll_seq[41]  `endif
                                        `ifdef STREAM41_OUT_WIDTH | stream_out_desc_poll_seq[41] `endif
                                        `ifdef STREAM42_IN_WIDTH  | stream_in_desc_poll_seq[42]  `endif
                                        `ifdef STREAM42_OUT_WIDTH | stream_out_desc_poll_seq[42] `endif
                                        `ifdef STREAM43_IN_WIDTH  | stream_in_desc_poll_seq[43]  `endif
                                        `ifdef STREAM43_OUT_WIDTH | stream_out_desc_poll_seq[43] `endif
                                        `ifdef STREAM44_IN_WIDTH  | stream_in_desc_poll_seq[44]  `endif
                                        `ifdef STREAM44_OUT_WIDTH | stream_out_desc_poll_seq[44] `endif
                                        `ifdef STREAM45_IN_WIDTH  | stream_in_desc_poll_seq[45]  `endif
                                        `ifdef STREAM45_OUT_WIDTH | stream_out_desc_poll_seq[45] `endif
                                        `ifdef STREAM46_IN_WIDTH  | stream_in_desc_poll_seq[46]  `endif
                                        `ifdef STREAM46_OUT_WIDTH | stream_out_desc_poll_seq[46] `endif
                                        `ifdef STREAM47_IN_WIDTH  | stream_in_desc_poll_seq[47]  `endif
                                        `ifdef STREAM47_OUT_WIDTH | stream_out_desc_poll_seq[47] `endif
                                        `ifdef STREAM48_IN_WIDTH  | stream_in_desc_poll_seq[48]  `endif
                                        `ifdef STREAM48_OUT_WIDTH | stream_out_desc_poll_seq[48] `endif
                                        `ifdef STREAM49_IN_WIDTH  | stream_in_desc_poll_seq[49]  `endif
                                        `ifdef STREAM49_OUT_WIDTH | stream_out_desc_poll_seq[49] `endif
                                        `ifdef STREAM50_IN_WIDTH  | stream_in_desc_poll_seq[50]  `endif
                                        `ifdef STREAM50_OUT_WIDTH | stream_out_desc_poll_seq[50] `endif
                                        `ifdef STREAM51_IN_WIDTH  | stream_in_desc_poll_seq[51]  `endif
                                        `ifdef STREAM51_OUT_WIDTH | stream_out_desc_poll_seq[51] `endif
                                        `ifdef STREAM52_IN_WIDTH  | stream_in_desc_poll_seq[52]  `endif
                                        `ifdef STREAM52_OUT_WIDTH | stream_out_desc_poll_seq[52] `endif
                                        `ifdef STREAM53_IN_WIDTH  | stream_in_desc_poll_seq[53]  `endif
                                        `ifdef STREAM53_OUT_WIDTH | stream_out_desc_poll_seq[53] `endif
                                        `ifdef STREAM54_IN_WIDTH  | stream_in_desc_poll_seq[54]  `endif
                                        `ifdef STREAM54_OUT_WIDTH | stream_out_desc_poll_seq[54] `endif
                                        `ifdef STREAM55_IN_WIDTH  | stream_in_desc_poll_seq[55]  `endif
                                        `ifdef STREAM55_OUT_WIDTH | stream_out_desc_poll_seq[55] `endif
                                        `ifdef STREAM56_IN_WIDTH  | stream_in_desc_poll_seq[56]  `endif
                                        `ifdef STREAM56_OUT_WIDTH | stream_out_desc_poll_seq[56] `endif
                                        `ifdef STREAM57_IN_WIDTH  | stream_in_desc_poll_seq[57]  `endif
                                        `ifdef STREAM57_OUT_WIDTH | stream_out_desc_poll_seq[57] `endif
                                        `ifdef STREAM58_IN_WIDTH  | stream_in_desc_poll_seq[58]  `endif
                                        `ifdef STREAM58_OUT_WIDTH | stream_out_desc_poll_seq[58] `endif
                                        `ifdef STREAM59_IN_WIDTH  | stream_in_desc_poll_seq[59]  `endif
                                        `ifdef STREAM59_OUT_WIDTH | stream_out_desc_poll_seq[59] `endif
                                        `ifdef STREAM60_IN_WIDTH  | stream_in_desc_poll_seq[60]  `endif
                                        `ifdef STREAM60_OUT_WIDTH | stream_out_desc_poll_seq[60] `endif
                                        `ifdef STREAM61_IN_WIDTH  | stream_in_desc_poll_seq[61]  `endif
                                        `ifdef STREAM61_OUT_WIDTH | stream_out_desc_poll_seq[61] `endif
                                        `ifdef STREAM62_IN_WIDTH  | stream_in_desc_poll_seq[62]  `endif
                                        `ifdef STREAM62_OUT_WIDTH | stream_out_desc_poll_seq[62] `endif
                                        `ifdef STREAM63_IN_WIDTH  | stream_in_desc_poll_seq[63]  `endif
                                        `ifdef STREAM63_OUT_WIDTH | stream_out_desc_poll_seq[63] `endif
                                        `ifdef STREAM64_IN_WIDTH  | stream_in_desc_poll_seq[64]  `endif
                                        `ifdef STREAM64_OUT_WIDTH | stream_out_desc_poll_seq[64] `endif
                                        `ifdef STREAM65_IN_WIDTH  | stream_in_desc_poll_seq[65]  `endif
                                        `ifdef STREAM65_OUT_WIDTH | stream_out_desc_poll_seq[65] `endif
                                        `ifdef STREAM66_IN_WIDTH  | stream_in_desc_poll_seq[66]  `endif
                                        `ifdef STREAM66_OUT_WIDTH | stream_out_desc_poll_seq[66] `endif
                                        `ifdef STREAM67_IN_WIDTH  | stream_in_desc_poll_seq[67]  `endif
                                        `ifdef STREAM67_OUT_WIDTH | stream_out_desc_poll_seq[67] `endif
                                        `ifdef STREAM68_IN_WIDTH  | stream_in_desc_poll_seq[68]  `endif
                                        `ifdef STREAM68_OUT_WIDTH | stream_out_desc_poll_seq[68] `endif
                                        `ifdef STREAM69_IN_WIDTH  | stream_in_desc_poll_seq[69]  `endif
                                        `ifdef STREAM69_OUT_WIDTH | stream_out_desc_poll_seq[69] `endif
                                        `ifdef STREAM70_IN_WIDTH  | stream_in_desc_poll_seq[70]  `endif
                                        `ifdef STREAM70_OUT_WIDTH | stream_out_desc_poll_seq[70] `endif
                                        `ifdef STREAM71_IN_WIDTH  | stream_in_desc_poll_seq[71]  `endif
                                        `ifdef STREAM71_OUT_WIDTH | stream_out_desc_poll_seq[71] `endif
                                        `ifdef STREAM72_IN_WIDTH  | stream_in_desc_poll_seq[72]  `endif
                                        `ifdef STREAM72_OUT_WIDTH | stream_out_desc_poll_seq[72] `endif
                                        `ifdef STREAM73_IN_WIDTH  | stream_in_desc_poll_seq[73]  `endif
                                        `ifdef STREAM73_OUT_WIDTH | stream_out_desc_poll_seq[73] `endif
                                        `ifdef STREAM74_IN_WIDTH  | stream_in_desc_poll_seq[74]  `endif
                                        `ifdef STREAM74_OUT_WIDTH | stream_out_desc_poll_seq[74] `endif
                                        `ifdef STREAM75_IN_WIDTH  | stream_in_desc_poll_seq[75]  `endif
                                        `ifdef STREAM75_OUT_WIDTH | stream_out_desc_poll_seq[75] `endif
                                        `ifdef STREAM76_IN_WIDTH  | stream_in_desc_poll_seq[76]  `endif
                                        `ifdef STREAM76_OUT_WIDTH | stream_out_desc_poll_seq[76] `endif
                                        `ifdef STREAM77_IN_WIDTH  | stream_in_desc_poll_seq[77]  `endif
                                        `ifdef STREAM77_OUT_WIDTH | stream_out_desc_poll_seq[77] `endif
                                        `ifdef STREAM78_IN_WIDTH  | stream_in_desc_poll_seq[78]  `endif
                                        `ifdef STREAM78_OUT_WIDTH | stream_out_desc_poll_seq[78] `endif
                                        `ifdef STREAM79_IN_WIDTH  | stream_in_desc_poll_seq[79]  `endif
                                        `ifdef STREAM79_OUT_WIDTH | stream_out_desc_poll_seq[79] `endif
                                        `ifdef STREAM80_IN_WIDTH  | stream_in_desc_poll_seq[80]  `endif
                                        `ifdef STREAM80_OUT_WIDTH | stream_out_desc_poll_seq[80] `endif
                                        `ifdef STREAM81_IN_WIDTH  | stream_in_desc_poll_seq[81]  `endif
                                        `ifdef STREAM81_OUT_WIDTH | stream_out_desc_poll_seq[81] `endif
                                        `ifdef STREAM82_IN_WIDTH  | stream_in_desc_poll_seq[82]  `endif
                                        `ifdef STREAM82_OUT_WIDTH | stream_out_desc_poll_seq[82] `endif
                                        `ifdef STREAM83_IN_WIDTH  | stream_in_desc_poll_seq[83]  `endif
                                        `ifdef STREAM83_OUT_WIDTH | stream_out_desc_poll_seq[83] `endif
                                        `ifdef STREAM84_IN_WIDTH  | stream_in_desc_poll_seq[84]  `endif
                                        `ifdef STREAM84_OUT_WIDTH | stream_out_desc_poll_seq[84] `endif
                                        `ifdef STREAM85_IN_WIDTH  | stream_in_desc_poll_seq[85]  `endif
                                        `ifdef STREAM85_OUT_WIDTH | stream_out_desc_poll_seq[85] `endif
                                        `ifdef STREAM86_IN_WIDTH  | stream_in_desc_poll_seq[86]  `endif
                                        `ifdef STREAM86_OUT_WIDTH | stream_out_desc_poll_seq[86] `endif
                                        `ifdef STREAM87_IN_WIDTH  | stream_in_desc_poll_seq[87]  `endif
                                        `ifdef STREAM87_OUT_WIDTH | stream_out_desc_poll_seq[87] `endif
                                        `ifdef STREAM88_IN_WIDTH  | stream_in_desc_poll_seq[88]  `endif
                                        `ifdef STREAM88_OUT_WIDTH | stream_out_desc_poll_seq[88] `endif
                                        `ifdef STREAM89_IN_WIDTH  | stream_in_desc_poll_seq[89]  `endif
                                        `ifdef STREAM89_OUT_WIDTH | stream_out_desc_poll_seq[89] `endif
                                        `ifdef STREAM90_IN_WIDTH  | stream_in_desc_poll_seq[90]  `endif
                                        `ifdef STREAM90_OUT_WIDTH | stream_out_desc_poll_seq[90] `endif
                                        `ifdef STREAM91_IN_WIDTH  | stream_in_desc_poll_seq[91]  `endif
                                        `ifdef STREAM91_OUT_WIDTH | stream_out_desc_poll_seq[91] `endif
                                        `ifdef STREAM92_IN_WIDTH  | stream_in_desc_poll_seq[92]  `endif
                                        `ifdef STREAM92_OUT_WIDTH | stream_out_desc_poll_seq[92] `endif
                                        `ifdef STREAM93_IN_WIDTH  | stream_in_desc_poll_seq[93]  `endif
                                        `ifdef STREAM93_OUT_WIDTH | stream_out_desc_poll_seq[93] `endif
                                        `ifdef STREAM94_IN_WIDTH  | stream_in_desc_poll_seq[94]  `endif
                                        `ifdef STREAM94_OUT_WIDTH | stream_out_desc_poll_seq[94] `endif
                                        `ifdef STREAM95_IN_WIDTH  | stream_in_desc_poll_seq[95]  `endif
                                        `ifdef STREAM95_OUT_WIDTH | stream_out_desc_poll_seq[95] `endif
                                        `ifdef STREAM96_IN_WIDTH  | stream_in_desc_poll_seq[96]  `endif
                                        `ifdef STREAM96_OUT_WIDTH | stream_out_desc_poll_seq[96] `endif
                                        `ifdef STREAM97_IN_WIDTH  | stream_in_desc_poll_seq[97]  `endif
                                        `ifdef STREAM97_OUT_WIDTH | stream_out_desc_poll_seq[97] `endif
                                        `ifdef STREAM98_IN_WIDTH  | stream_in_desc_poll_seq[98]  `endif
                                        `ifdef STREAM98_OUT_WIDTH | stream_out_desc_poll_seq[98] `endif
                                        `ifdef STREAM99_IN_WIDTH  | stream_in_desc_poll_seq[99]  `endif
                                        `ifdef STREAM99_OUT_WIDTH | stream_out_desc_poll_seq[99] `endif
                                        `ifdef STREAM100_IN_WIDTH  | stream_in_desc_poll_seq[100]  `endif
                                        `ifdef STREAM100_OUT_WIDTH | stream_out_desc_poll_seq[100] `endif
                                        `ifdef STREAM101_IN_WIDTH  | stream_in_desc_poll_seq[101]  `endif
                                        `ifdef STREAM101_OUT_WIDTH | stream_out_desc_poll_seq[101] `endif
                                        `ifdef STREAM102_IN_WIDTH  | stream_in_desc_poll_seq[102]  `endif
                                        `ifdef STREAM102_OUT_WIDTH | stream_out_desc_poll_seq[102] `endif
                                        `ifdef STREAM103_IN_WIDTH  | stream_in_desc_poll_seq[103]  `endif
                                        `ifdef STREAM103_OUT_WIDTH | stream_out_desc_poll_seq[103] `endif
                                        `ifdef STREAM104_IN_WIDTH  | stream_in_desc_poll_seq[104]  `endif
                                        `ifdef STREAM104_OUT_WIDTH | stream_out_desc_poll_seq[104] `endif
                                        `ifdef STREAM105_IN_WIDTH  | stream_in_desc_poll_seq[105]  `endif
                                        `ifdef STREAM105_OUT_WIDTH | stream_out_desc_poll_seq[105] `endif
                                        `ifdef STREAM106_IN_WIDTH  | stream_in_desc_poll_seq[106]  `endif
                                        `ifdef STREAM106_OUT_WIDTH | stream_out_desc_poll_seq[106] `endif
                                        `ifdef STREAM107_IN_WIDTH  | stream_in_desc_poll_seq[107]  `endif
                                        `ifdef STREAM107_OUT_WIDTH | stream_out_desc_poll_seq[107] `endif
                                        `ifdef STREAM108_IN_WIDTH  | stream_in_desc_poll_seq[108]  `endif
                                        `ifdef STREAM108_OUT_WIDTH | stream_out_desc_poll_seq[108] `endif
                                        `ifdef STREAM109_IN_WIDTH  | stream_in_desc_poll_seq[109]  `endif
                                        `ifdef STREAM109_OUT_WIDTH | stream_out_desc_poll_seq[109] `endif
                                        `ifdef STREAM110_IN_WIDTH  | stream_in_desc_poll_seq[110]  `endif
                                        `ifdef STREAM110_OUT_WIDTH | stream_out_desc_poll_seq[110] `endif
                                        `ifdef STREAM111_IN_WIDTH  | stream_in_desc_poll_seq[111]  `endif
                                        `ifdef STREAM111_OUT_WIDTH | stream_out_desc_poll_seq[111] `endif
                                        `ifdef STREAM112_IN_WIDTH  | stream_in_desc_poll_seq[112]  `endif
                                        `ifdef STREAM112_OUT_WIDTH | stream_out_desc_poll_seq[112] `endif
                                        `ifdef STREAM113_IN_WIDTH  | stream_in_desc_poll_seq[113]  `endif
                                        `ifdef STREAM113_OUT_WIDTH | stream_out_desc_poll_seq[113] `endif
                                        `ifdef STREAM114_IN_WIDTH  | stream_in_desc_poll_seq[114]  `endif
                                        `ifdef STREAM114_OUT_WIDTH | stream_out_desc_poll_seq[114] `endif
                                        `ifdef STREAM115_IN_WIDTH  | stream_in_desc_poll_seq[115]  `endif
                                        `ifdef STREAM115_OUT_WIDTH | stream_out_desc_poll_seq[115] `endif
                                        `ifdef STREAM116_IN_WIDTH  | stream_in_desc_poll_seq[116]  `endif
                                        `ifdef STREAM116_OUT_WIDTH | stream_out_desc_poll_seq[116] `endif
                                        `ifdef STREAM117_IN_WIDTH  | stream_in_desc_poll_seq[117]  `endif
                                        `ifdef STREAM117_OUT_WIDTH | stream_out_desc_poll_seq[117] `endif
                                        `ifdef STREAM118_IN_WIDTH  | stream_in_desc_poll_seq[118]  `endif
                                        `ifdef STREAM118_OUT_WIDTH | stream_out_desc_poll_seq[118] `endif
                                        `ifdef STREAM119_IN_WIDTH  | stream_in_desc_poll_seq[119]  `endif
                                        `ifdef STREAM119_OUT_WIDTH | stream_out_desc_poll_seq[119] `endif
                                        `ifdef STREAM120_IN_WIDTH  | stream_in_desc_poll_seq[120]  `endif
                                        `ifdef STREAM120_OUT_WIDTH | stream_out_desc_poll_seq[120] `endif
                                        `ifdef STREAM121_IN_WIDTH  | stream_in_desc_poll_seq[121]  `endif
                                        `ifdef STREAM121_OUT_WIDTH | stream_out_desc_poll_seq[121] `endif
                                        `ifdef STREAM122_IN_WIDTH  | stream_in_desc_poll_seq[122]  `endif
                                        `ifdef STREAM122_OUT_WIDTH | stream_out_desc_poll_seq[122] `endif
                                        `ifdef STREAM123_IN_WIDTH  | stream_in_desc_poll_seq[123]  `endif
                                        `ifdef STREAM123_OUT_WIDTH | stream_out_desc_poll_seq[123] `endif
                                        `ifdef STREAM124_IN_WIDTH  | stream_in_desc_poll_seq[124]  `endif
                                        `ifdef STREAM124_OUT_WIDTH | stream_out_desc_poll_seq[124] `endif
                                        `ifdef STREAM125_IN_WIDTH  | stream_in_desc_poll_seq[125]  `endif
                                        `ifdef STREAM125_OUT_WIDTH | stream_out_desc_poll_seq[125] `endif
                                        `ifdef STREAM126_IN_WIDTH  | stream_in_desc_poll_seq[126]  `endif
                                        `ifdef STREAM126_OUT_WIDTH | stream_out_desc_poll_seq[126] `endif
                                        );
    assign s_poll_next_desc_valid   = (1'b0
                                        `ifdef PICOBUS_WIDTH  | s_poll_next_desc_valid_userpb `endif
                                        `ifdef STREAM1_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[1]  `endif
                                        `ifdef STREAM1_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[1] `endif
                                        `ifdef STREAM2_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[2]  `endif
                                        `ifdef STREAM2_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[2] `endif
                                        `ifdef STREAM3_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[3]  `endif
                                        `ifdef STREAM3_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[3] `endif
                                        `ifdef STREAM4_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[4]  `endif
                                        `ifdef STREAM4_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[4] `endif
                                        `ifdef STREAM5_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[5]  `endif
                                        `ifdef STREAM5_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[5] `endif
                                        `ifdef STREAM6_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[6]  `endif
                                        `ifdef STREAM6_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[6] `endif
                                        `ifdef STREAM7_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[7]  `endif
                                        `ifdef STREAM7_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[7] `endif
                                        `ifdef STREAM8_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[8]  `endif
                                        `ifdef STREAM8_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[8] `endif
                                        `ifdef STREAM9_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[9]  `endif
                                        `ifdef STREAM9_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[9] `endif
                                        `ifdef STREAM10_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[10]  `endif
                                        `ifdef STREAM10_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[10] `endif
                                        `ifdef STREAM11_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[11]  `endif
                                        `ifdef STREAM11_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[11] `endif
                                        `ifdef STREAM12_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[12]  `endif
                                        `ifdef STREAM12_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[12] `endif
                                        `ifdef STREAM13_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[13]  `endif
                                        `ifdef STREAM13_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[13] `endif
                                        `ifdef STREAM14_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[14]  `endif
                                        `ifdef STREAM14_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[14] `endif
                                        `ifdef STREAM15_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[15]  `endif
                                        `ifdef STREAM15_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[15] `endif
                                        `ifdef STREAM16_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[16]  `endif
                                        `ifdef STREAM16_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[16] `endif
                                        `ifdef STREAM17_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[17]  `endif
                                        `ifdef STREAM17_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[17] `endif
                                        `ifdef STREAM18_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[18]  `endif
                                        `ifdef STREAM18_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[18] `endif
                                        `ifdef STREAM19_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[19]  `endif
                                        `ifdef STREAM19_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[19] `endif
                                        `ifdef STREAM20_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[20]  `endif
                                        `ifdef STREAM20_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[20] `endif
                                        `ifdef STREAM21_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[21]  `endif
                                        `ifdef STREAM21_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[21] `endif
                                        `ifdef STREAM22_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[22]  `endif
                                        `ifdef STREAM22_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[22] `endif
                                        `ifdef STREAM23_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[23]  `endif
                                        `ifdef STREAM23_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[23] `endif
                                        `ifdef STREAM24_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[24]  `endif
                                        `ifdef STREAM24_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[24] `endif
                                        `ifdef STREAM25_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[25]  `endif
                                        `ifdef STREAM25_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[25] `endif
                                        `ifdef STREAM26_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[26]  `endif
                                        `ifdef STREAM26_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[26] `endif
                                        `ifdef STREAM27_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[27]  `endif
                                        `ifdef STREAM27_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[27] `endif
                                        `ifdef STREAM28_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[28]  `endif
                                        `ifdef STREAM28_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[28] `endif
                                        `ifdef STREAM29_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[29]  `endif
                                        `ifdef STREAM29_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[29] `endif
                                        `ifdef STREAM30_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[30]  `endif
                                        `ifdef STREAM30_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[30] `endif
                                        `ifdef STREAM31_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[31]  `endif
                                        `ifdef STREAM31_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[31] `endif
                                        `ifdef STREAM32_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[32]  `endif
                                        `ifdef STREAM32_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[32] `endif
                                        `ifdef STREAM33_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[33]  `endif
                                        `ifdef STREAM33_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[33] `endif
                                        `ifdef STREAM34_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[34]  `endif
                                        `ifdef STREAM34_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[34] `endif
                                        `ifdef STREAM35_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[35]  `endif
                                        `ifdef STREAM35_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[35] `endif
                                        `ifdef STREAM36_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[36]  `endif
                                        `ifdef STREAM36_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[36] `endif
                                        `ifdef STREAM37_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[37]  `endif
                                        `ifdef STREAM37_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[37] `endif
                                        `ifdef STREAM38_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[38]  `endif
                                        `ifdef STREAM38_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[38] `endif
                                        `ifdef STREAM39_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[39]  `endif
                                        `ifdef STREAM39_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[39] `endif
                                        `ifdef STREAM40_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[40]  `endif
                                        `ifdef STREAM40_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[40] `endif
                                        `ifdef STREAM41_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[41]  `endif
                                        `ifdef STREAM41_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[41] `endif
                                        `ifdef STREAM42_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[42]  `endif
                                        `ifdef STREAM42_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[42] `endif
                                        `ifdef STREAM43_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[43]  `endif
                                        `ifdef STREAM43_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[43] `endif
                                        `ifdef STREAM44_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[44]  `endif
                                        `ifdef STREAM44_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[44] `endif
                                        `ifdef STREAM45_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[45]  `endif
                                        `ifdef STREAM45_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[45] `endif
                                        `ifdef STREAM46_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[46]  `endif
                                        `ifdef STREAM46_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[46] `endif
                                        `ifdef STREAM47_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[47]  `endif
                                        `ifdef STREAM47_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[47] `endif
                                        `ifdef STREAM48_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[48]  `endif
                                        `ifdef STREAM48_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[48] `endif
                                        `ifdef STREAM49_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[49]  `endif
                                        `ifdef STREAM49_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[49] `endif
                                        `ifdef STREAM50_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[50]  `endif
                                        `ifdef STREAM50_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[50] `endif
                                        `ifdef STREAM51_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[51]  `endif
                                        `ifdef STREAM51_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[51] `endif
                                        `ifdef STREAM52_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[52]  `endif
                                        `ifdef STREAM52_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[52] `endif
                                        `ifdef STREAM53_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[53]  `endif
                                        `ifdef STREAM53_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[53] `endif
                                        `ifdef STREAM54_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[54]  `endif
                                        `ifdef STREAM54_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[54] `endif
                                        `ifdef STREAM55_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[55]  `endif
                                        `ifdef STREAM55_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[55] `endif
                                        `ifdef STREAM56_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[56]  `endif
                                        `ifdef STREAM56_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[56] `endif
                                        `ifdef STREAM57_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[57]  `endif
                                        `ifdef STREAM57_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[57] `endif
                                        `ifdef STREAM58_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[58]  `endif
                                        `ifdef STREAM58_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[58] `endif
                                        `ifdef STREAM59_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[59]  `endif
                                        `ifdef STREAM59_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[59] `endif
                                        `ifdef STREAM60_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[60]  `endif
                                        `ifdef STREAM60_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[60] `endif
                                        `ifdef STREAM61_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[61]  `endif
                                        `ifdef STREAM61_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[61] `endif
                                        `ifdef STREAM62_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[62]  `endif
                                        `ifdef STREAM62_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[62] `endif
                                        `ifdef STREAM63_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[63]  `endif
                                        `ifdef STREAM63_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[63] `endif
                                        `ifdef STREAM64_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[64]  `endif
                                        `ifdef STREAM64_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[64] `endif
                                        `ifdef STREAM65_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[65]  `endif
                                        `ifdef STREAM65_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[65] `endif
                                        `ifdef STREAM66_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[66]  `endif
                                        `ifdef STREAM66_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[66] `endif
                                        `ifdef STREAM67_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[67]  `endif
                                        `ifdef STREAM67_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[67] `endif
                                        `ifdef STREAM68_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[68]  `endif
                                        `ifdef STREAM68_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[68] `endif
                                        `ifdef STREAM69_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[69]  `endif
                                        `ifdef STREAM69_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[69] `endif
                                        `ifdef STREAM70_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[70]  `endif
                                        `ifdef STREAM70_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[70] `endif
                                        `ifdef STREAM71_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[71]  `endif
                                        `ifdef STREAM71_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[71] `endif
                                        `ifdef STREAM72_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[72]  `endif
                                        `ifdef STREAM72_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[72] `endif
                                        `ifdef STREAM73_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[73]  `endif
                                        `ifdef STREAM73_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[73] `endif
                                        `ifdef STREAM74_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[74]  `endif
                                        `ifdef STREAM74_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[74] `endif
                                        `ifdef STREAM75_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[75]  `endif
                                        `ifdef STREAM75_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[75] `endif
                                        `ifdef STREAM76_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[76]  `endif
                                        `ifdef STREAM76_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[76] `endif
                                        `ifdef STREAM77_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[77]  `endif
                                        `ifdef STREAM77_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[77] `endif
                                        `ifdef STREAM78_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[78]  `endif
                                        `ifdef STREAM78_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[78] `endif
                                        `ifdef STREAM79_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[79]  `endif
                                        `ifdef STREAM79_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[79] `endif
                                        `ifdef STREAM80_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[80]  `endif
                                        `ifdef STREAM80_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[80] `endif
                                        `ifdef STREAM81_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[81]  `endif
                                        `ifdef STREAM81_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[81] `endif
                                        `ifdef STREAM82_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[82]  `endif
                                        `ifdef STREAM82_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[82] `endif
                                        `ifdef STREAM83_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[83]  `endif
                                        `ifdef STREAM83_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[83] `endif
                                        `ifdef STREAM84_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[84]  `endif
                                        `ifdef STREAM84_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[84] `endif
                                        `ifdef STREAM85_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[85]  `endif
                                        `ifdef STREAM85_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[85] `endif
                                        `ifdef STREAM86_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[86]  `endif
                                        `ifdef STREAM86_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[86] `endif
                                        `ifdef STREAM87_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[87]  `endif
                                        `ifdef STREAM87_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[87] `endif
                                        `ifdef STREAM88_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[88]  `endif
                                        `ifdef STREAM88_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[88] `endif
                                        `ifdef STREAM89_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[89]  `endif
                                        `ifdef STREAM89_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[89] `endif
                                        `ifdef STREAM90_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[90]  `endif
                                        `ifdef STREAM90_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[90] `endif
                                        `ifdef STREAM91_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[91]  `endif
                                        `ifdef STREAM91_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[91] `endif
                                        `ifdef STREAM92_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[92]  `endif
                                        `ifdef STREAM92_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[92] `endif
                                        `ifdef STREAM93_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[93]  `endif
                                        `ifdef STREAM93_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[93] `endif
                                        `ifdef STREAM94_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[94]  `endif
                                        `ifdef STREAM94_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[94] `endif
                                        `ifdef STREAM95_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[95]  `endif
                                        `ifdef STREAM95_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[95] `endif
                                        `ifdef STREAM96_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[96]  `endif
                                        `ifdef STREAM96_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[96] `endif
                                        `ifdef STREAM97_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[97]  `endif
                                        `ifdef STREAM97_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[97] `endif
                                        `ifdef STREAM98_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[98]  `endif
                                        `ifdef STREAM98_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[98] `endif
                                        `ifdef STREAM99_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[99]  `endif
                                        `ifdef STREAM99_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[99] `endif
                                        `ifdef STREAM100_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[100]  `endif
                                        `ifdef STREAM100_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[100] `endif
                                        `ifdef STREAM101_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[101]  `endif
                                        `ifdef STREAM101_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[101] `endif
                                        `ifdef STREAM102_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[102]  `endif
                                        `ifdef STREAM102_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[102] `endif
                                        `ifdef STREAM103_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[103]  `endif
                                        `ifdef STREAM103_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[103] `endif
                                        `ifdef STREAM104_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[104]  `endif
                                        `ifdef STREAM104_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[104] `endif
                                        `ifdef STREAM105_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[105]  `endif
                                        `ifdef STREAM105_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[105] `endif
                                        `ifdef STREAM106_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[106]  `endif
                                        `ifdef STREAM106_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[106] `endif
                                        `ifdef STREAM107_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[107]  `endif
                                        `ifdef STREAM107_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[107] `endif
                                        `ifdef STREAM108_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[108]  `endif
                                        `ifdef STREAM108_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[108] `endif
                                        `ifdef STREAM109_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[109]  `endif
                                        `ifdef STREAM109_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[109] `endif
                                        `ifdef STREAM110_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[110]  `endif
                                        `ifdef STREAM110_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[110] `endif
                                        `ifdef STREAM111_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[111]  `endif
                                        `ifdef STREAM111_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[111] `endif
                                        `ifdef STREAM112_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[112]  `endif
                                        `ifdef STREAM112_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[112] `endif
                                        `ifdef STREAM113_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[113]  `endif
                                        `ifdef STREAM113_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[113] `endif
                                        `ifdef STREAM114_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[114]  `endif
                                        `ifdef STREAM114_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[114] `endif
                                        `ifdef STREAM115_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[115]  `endif
                                        `ifdef STREAM115_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[115] `endif
                                        `ifdef STREAM116_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[116]  `endif
                                        `ifdef STREAM116_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[116] `endif
                                        `ifdef STREAM117_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[117]  `endif
                                        `ifdef STREAM117_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[117] `endif
                                        `ifdef STREAM118_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[118]  `endif
                                        `ifdef STREAM118_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[118] `endif
                                        `ifdef STREAM119_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[119]  `endif
                                        `ifdef STREAM119_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[119] `endif
                                        `ifdef STREAM120_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[120]  `endif
                                        `ifdef STREAM120_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[120] `endif
                                        `ifdef STREAM121_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[121]  `endif
                                        `ifdef STREAM121_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[121] `endif
                                        `ifdef STREAM122_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[122]  `endif
                                        `ifdef STREAM122_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[122] `endif
                                        `ifdef STREAM123_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[123]  `endif
                                        `ifdef STREAM123_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[123] `endif
                                        `ifdef STREAM124_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[124]  `endif
                                        `ifdef STREAM124_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[124] `endif
                                        `ifdef STREAM125_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[125]  `endif
                                        `ifdef STREAM125_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[125] `endif
                                        `ifdef STREAM126_IN_WIDTH  | stream_in_desc_poll_next_desc_valid[126]  `endif
                                        `ifdef STREAM126_OUT_WIDTH | stream_out_desc_poll_next_desc_valid[126] `endif
                                        );
    assign s_poll_next_desc[127:0]  = (128'h0
                                        `ifdef PICOBUS_WIDTH | s_poll_next_desc_userpb    `endif
                                        `ifdef STREAM1_IN_WIDTH  | stream_in_desc_poll_next_desc[1]  `endif
                                        `ifdef STREAM1_OUT_WIDTH | stream_out_desc_poll_next_desc[1] `endif
                                        `ifdef STREAM2_IN_WIDTH  | stream_in_desc_poll_next_desc[2]  `endif
                                        `ifdef STREAM2_OUT_WIDTH | stream_out_desc_poll_next_desc[2] `endif
                                        `ifdef STREAM3_IN_WIDTH  | stream_in_desc_poll_next_desc[3]  `endif
                                        `ifdef STREAM3_OUT_WIDTH | stream_out_desc_poll_next_desc[3] `endif
                                        `ifdef STREAM4_IN_WIDTH  | stream_in_desc_poll_next_desc[4]  `endif
                                        `ifdef STREAM4_OUT_WIDTH | stream_out_desc_poll_next_desc[4] `endif
                                        `ifdef STREAM5_IN_WIDTH  | stream_in_desc_poll_next_desc[5]  `endif
                                        `ifdef STREAM5_OUT_WIDTH | stream_out_desc_poll_next_desc[5] `endif
                                        `ifdef STREAM6_IN_WIDTH  | stream_in_desc_poll_next_desc[6]  `endif
                                        `ifdef STREAM6_OUT_WIDTH | stream_out_desc_poll_next_desc[6] `endif
                                        `ifdef STREAM7_IN_WIDTH  | stream_in_desc_poll_next_desc[7]  `endif
                                        `ifdef STREAM7_OUT_WIDTH | stream_out_desc_poll_next_desc[7] `endif
                                        `ifdef STREAM8_IN_WIDTH  | stream_in_desc_poll_next_desc[8]  `endif
                                        `ifdef STREAM8_OUT_WIDTH | stream_out_desc_poll_next_desc[8] `endif
                                        `ifdef STREAM9_IN_WIDTH  | stream_in_desc_poll_next_desc[9]  `endif
                                        `ifdef STREAM9_OUT_WIDTH | stream_out_desc_poll_next_desc[9] `endif
                                        `ifdef STREAM10_IN_WIDTH  | stream_in_desc_poll_next_desc[10]  `endif
                                        `ifdef STREAM10_OUT_WIDTH | stream_out_desc_poll_next_desc[10] `endif
                                        `ifdef STREAM11_IN_WIDTH  | stream_in_desc_poll_next_desc[11]  `endif
                                        `ifdef STREAM11_OUT_WIDTH | stream_out_desc_poll_next_desc[11] `endif
                                        `ifdef STREAM12_IN_WIDTH  | stream_in_desc_poll_next_desc[12]  `endif
                                        `ifdef STREAM12_OUT_WIDTH | stream_out_desc_poll_next_desc[12] `endif
                                        `ifdef STREAM13_IN_WIDTH  | stream_in_desc_poll_next_desc[13]  `endif
                                        `ifdef STREAM13_OUT_WIDTH | stream_out_desc_poll_next_desc[13] `endif
                                        `ifdef STREAM14_IN_WIDTH  | stream_in_desc_poll_next_desc[14]  `endif
                                        `ifdef STREAM14_OUT_WIDTH | stream_out_desc_poll_next_desc[14] `endif
                                        `ifdef STREAM15_IN_WIDTH  | stream_in_desc_poll_next_desc[15]  `endif
                                        `ifdef STREAM15_OUT_WIDTH | stream_out_desc_poll_next_desc[15] `endif
                                        `ifdef STREAM16_IN_WIDTH  | stream_in_desc_poll_next_desc[16]  `endif
                                        `ifdef STREAM16_OUT_WIDTH | stream_out_desc_poll_next_desc[16] `endif
                                        `ifdef STREAM17_IN_WIDTH  | stream_in_desc_poll_next_desc[17]  `endif
                                        `ifdef STREAM17_OUT_WIDTH | stream_out_desc_poll_next_desc[17] `endif
                                        `ifdef STREAM18_IN_WIDTH  | stream_in_desc_poll_next_desc[18]  `endif
                                        `ifdef STREAM18_OUT_WIDTH | stream_out_desc_poll_next_desc[18] `endif
                                        `ifdef STREAM19_IN_WIDTH  | stream_in_desc_poll_next_desc[19]  `endif
                                        `ifdef STREAM19_OUT_WIDTH | stream_out_desc_poll_next_desc[19] `endif
                                        `ifdef STREAM20_IN_WIDTH  | stream_in_desc_poll_next_desc[20]  `endif
                                        `ifdef STREAM20_OUT_WIDTH | stream_out_desc_poll_next_desc[20] `endif
                                        `ifdef STREAM21_IN_WIDTH  | stream_in_desc_poll_next_desc[21]  `endif
                                        `ifdef STREAM21_OUT_WIDTH | stream_out_desc_poll_next_desc[21] `endif
                                        `ifdef STREAM22_IN_WIDTH  | stream_in_desc_poll_next_desc[22]  `endif
                                        `ifdef STREAM22_OUT_WIDTH | stream_out_desc_poll_next_desc[22] `endif
                                        `ifdef STREAM23_IN_WIDTH  | stream_in_desc_poll_next_desc[23]  `endif
                                        `ifdef STREAM23_OUT_WIDTH | stream_out_desc_poll_next_desc[23] `endif
                                        `ifdef STREAM24_IN_WIDTH  | stream_in_desc_poll_next_desc[24]  `endif
                                        `ifdef STREAM24_OUT_WIDTH | stream_out_desc_poll_next_desc[24] `endif
                                        `ifdef STREAM25_IN_WIDTH  | stream_in_desc_poll_next_desc[25]  `endif
                                        `ifdef STREAM25_OUT_WIDTH | stream_out_desc_poll_next_desc[25] `endif
                                        `ifdef STREAM26_IN_WIDTH  | stream_in_desc_poll_next_desc[26]  `endif
                                        `ifdef STREAM26_OUT_WIDTH | stream_out_desc_poll_next_desc[26] `endif
                                        `ifdef STREAM27_IN_WIDTH  | stream_in_desc_poll_next_desc[27]  `endif
                                        `ifdef STREAM27_OUT_WIDTH | stream_out_desc_poll_next_desc[27] `endif
                                        `ifdef STREAM28_IN_WIDTH  | stream_in_desc_poll_next_desc[28]  `endif
                                        `ifdef STREAM28_OUT_WIDTH | stream_out_desc_poll_next_desc[28] `endif
                                        `ifdef STREAM29_IN_WIDTH  | stream_in_desc_poll_next_desc[29]  `endif
                                        `ifdef STREAM29_OUT_WIDTH | stream_out_desc_poll_next_desc[29] `endif
                                        `ifdef STREAM30_IN_WIDTH  | stream_in_desc_poll_next_desc[30]  `endif
                                        `ifdef STREAM30_OUT_WIDTH | stream_out_desc_poll_next_desc[30] `endif
                                        `ifdef STREAM31_IN_WIDTH  | stream_in_desc_poll_next_desc[31]  `endif
                                        `ifdef STREAM31_OUT_WIDTH | stream_out_desc_poll_next_desc[31] `endif
                                        `ifdef STREAM32_IN_WIDTH  | stream_in_desc_poll_next_desc[32]  `endif
                                        `ifdef STREAM32_OUT_WIDTH | stream_out_desc_poll_next_desc[32] `endif
                                        `ifdef STREAM33_IN_WIDTH  | stream_in_desc_poll_next_desc[33]  `endif
                                        `ifdef STREAM33_OUT_WIDTH | stream_out_desc_poll_next_desc[33] `endif
                                        `ifdef STREAM34_IN_WIDTH  | stream_in_desc_poll_next_desc[34]  `endif
                                        `ifdef STREAM34_OUT_WIDTH | stream_out_desc_poll_next_desc[34] `endif
                                        `ifdef STREAM35_IN_WIDTH  | stream_in_desc_poll_next_desc[35]  `endif
                                        `ifdef STREAM35_OUT_WIDTH | stream_out_desc_poll_next_desc[35] `endif
                                        `ifdef STREAM36_IN_WIDTH  | stream_in_desc_poll_next_desc[36]  `endif
                                        `ifdef STREAM36_OUT_WIDTH | stream_out_desc_poll_next_desc[36] `endif
                                        `ifdef STREAM37_IN_WIDTH  | stream_in_desc_poll_next_desc[37]  `endif
                                        `ifdef STREAM37_OUT_WIDTH | stream_out_desc_poll_next_desc[37] `endif
                                        `ifdef STREAM38_IN_WIDTH  | stream_in_desc_poll_next_desc[38]  `endif
                                        `ifdef STREAM38_OUT_WIDTH | stream_out_desc_poll_next_desc[38] `endif
                                        `ifdef STREAM39_IN_WIDTH  | stream_in_desc_poll_next_desc[39]  `endif
                                        `ifdef STREAM39_OUT_WIDTH | stream_out_desc_poll_next_desc[39] `endif
                                        `ifdef STREAM40_IN_WIDTH  | stream_in_desc_poll_next_desc[40]  `endif
                                        `ifdef STREAM40_OUT_WIDTH | stream_out_desc_poll_next_desc[40] `endif
                                        `ifdef STREAM41_IN_WIDTH  | stream_in_desc_poll_next_desc[41]  `endif
                                        `ifdef STREAM41_OUT_WIDTH | stream_out_desc_poll_next_desc[41] `endif
                                        `ifdef STREAM42_IN_WIDTH  | stream_in_desc_poll_next_desc[42]  `endif
                                        `ifdef STREAM42_OUT_WIDTH | stream_out_desc_poll_next_desc[42] `endif
                                        `ifdef STREAM43_IN_WIDTH  | stream_in_desc_poll_next_desc[43]  `endif
                                        `ifdef STREAM43_OUT_WIDTH | stream_out_desc_poll_next_desc[43] `endif
                                        `ifdef STREAM44_IN_WIDTH  | stream_in_desc_poll_next_desc[44]  `endif
                                        `ifdef STREAM44_OUT_WIDTH | stream_out_desc_poll_next_desc[44] `endif
                                        `ifdef STREAM45_IN_WIDTH  | stream_in_desc_poll_next_desc[45]  `endif
                                        `ifdef STREAM45_OUT_WIDTH | stream_out_desc_poll_next_desc[45] `endif
                                        `ifdef STREAM46_IN_WIDTH  | stream_in_desc_poll_next_desc[46]  `endif
                                        `ifdef STREAM46_OUT_WIDTH | stream_out_desc_poll_next_desc[46] `endif
                                        `ifdef STREAM47_IN_WIDTH  | stream_in_desc_poll_next_desc[47]  `endif
                                        `ifdef STREAM47_OUT_WIDTH | stream_out_desc_poll_next_desc[47] `endif
                                        `ifdef STREAM48_IN_WIDTH  | stream_in_desc_poll_next_desc[48]  `endif
                                        `ifdef STREAM48_OUT_WIDTH | stream_out_desc_poll_next_desc[48] `endif
                                        `ifdef STREAM49_IN_WIDTH  | stream_in_desc_poll_next_desc[49]  `endif
                                        `ifdef STREAM49_OUT_WIDTH | stream_out_desc_poll_next_desc[49] `endif
                                        `ifdef STREAM50_IN_WIDTH  | stream_in_desc_poll_next_desc[50]  `endif
                                        `ifdef STREAM50_OUT_WIDTH | stream_out_desc_poll_next_desc[50] `endif
                                        `ifdef STREAM51_IN_WIDTH  | stream_in_desc_poll_next_desc[51]  `endif
                                        `ifdef STREAM51_OUT_WIDTH | stream_out_desc_poll_next_desc[51] `endif
                                        `ifdef STREAM52_IN_WIDTH  | stream_in_desc_poll_next_desc[52]  `endif
                                        `ifdef STREAM52_OUT_WIDTH | stream_out_desc_poll_next_desc[52] `endif
                                        `ifdef STREAM53_IN_WIDTH  | stream_in_desc_poll_next_desc[53]  `endif
                                        `ifdef STREAM53_OUT_WIDTH | stream_out_desc_poll_next_desc[53] `endif
                                        `ifdef STREAM54_IN_WIDTH  | stream_in_desc_poll_next_desc[54]  `endif
                                        `ifdef STREAM54_OUT_WIDTH | stream_out_desc_poll_next_desc[54] `endif
                                        `ifdef STREAM55_IN_WIDTH  | stream_in_desc_poll_next_desc[55]  `endif
                                        `ifdef STREAM55_OUT_WIDTH | stream_out_desc_poll_next_desc[55] `endif
                                        `ifdef STREAM56_IN_WIDTH  | stream_in_desc_poll_next_desc[56]  `endif
                                        `ifdef STREAM56_OUT_WIDTH | stream_out_desc_poll_next_desc[56] `endif
                                        `ifdef STREAM57_IN_WIDTH  | stream_in_desc_poll_next_desc[57]  `endif
                                        `ifdef STREAM57_OUT_WIDTH | stream_out_desc_poll_next_desc[57] `endif
                                        `ifdef STREAM58_IN_WIDTH  | stream_in_desc_poll_next_desc[58]  `endif
                                        `ifdef STREAM58_OUT_WIDTH | stream_out_desc_poll_next_desc[58] `endif
                                        `ifdef STREAM59_IN_WIDTH  | stream_in_desc_poll_next_desc[59]  `endif
                                        `ifdef STREAM59_OUT_WIDTH | stream_out_desc_poll_next_desc[59] `endif
                                        `ifdef STREAM60_IN_WIDTH  | stream_in_desc_poll_next_desc[60]  `endif
                                        `ifdef STREAM60_OUT_WIDTH | stream_out_desc_poll_next_desc[60] `endif
                                        `ifdef STREAM61_IN_WIDTH  | stream_in_desc_poll_next_desc[61]  `endif
                                        `ifdef STREAM61_OUT_WIDTH | stream_out_desc_poll_next_desc[61] `endif
                                        `ifdef STREAM62_IN_WIDTH  | stream_in_desc_poll_next_desc[62]  `endif
                                        `ifdef STREAM62_OUT_WIDTH | stream_out_desc_poll_next_desc[62] `endif
                                        `ifdef STREAM63_IN_WIDTH  | stream_in_desc_poll_next_desc[63]  `endif
                                        `ifdef STREAM63_OUT_WIDTH | stream_out_desc_poll_next_desc[63] `endif
                                        `ifdef STREAM64_IN_WIDTH  | stream_in_desc_poll_next_desc[64]  `endif
                                        `ifdef STREAM64_OUT_WIDTH | stream_out_desc_poll_next_desc[64] `endif
                                        `ifdef STREAM65_IN_WIDTH  | stream_in_desc_poll_next_desc[65]  `endif
                                        `ifdef STREAM65_OUT_WIDTH | stream_out_desc_poll_next_desc[65] `endif
                                        `ifdef STREAM66_IN_WIDTH  | stream_in_desc_poll_next_desc[66]  `endif
                                        `ifdef STREAM66_OUT_WIDTH | stream_out_desc_poll_next_desc[66] `endif
                                        `ifdef STREAM67_IN_WIDTH  | stream_in_desc_poll_next_desc[67]  `endif
                                        `ifdef STREAM67_OUT_WIDTH | stream_out_desc_poll_next_desc[67] `endif
                                        `ifdef STREAM68_IN_WIDTH  | stream_in_desc_poll_next_desc[68]  `endif
                                        `ifdef STREAM68_OUT_WIDTH | stream_out_desc_poll_next_desc[68] `endif
                                        `ifdef STREAM69_IN_WIDTH  | stream_in_desc_poll_next_desc[69]  `endif
                                        `ifdef STREAM69_OUT_WIDTH | stream_out_desc_poll_next_desc[69] `endif
                                        `ifdef STREAM70_IN_WIDTH  | stream_in_desc_poll_next_desc[70]  `endif
                                        `ifdef STREAM70_OUT_WIDTH | stream_out_desc_poll_next_desc[70] `endif
                                        `ifdef STREAM71_IN_WIDTH  | stream_in_desc_poll_next_desc[71]  `endif
                                        `ifdef STREAM71_OUT_WIDTH | stream_out_desc_poll_next_desc[71] `endif
                                        `ifdef STREAM72_IN_WIDTH  | stream_in_desc_poll_next_desc[72]  `endif
                                        `ifdef STREAM72_OUT_WIDTH | stream_out_desc_poll_next_desc[72] `endif
                                        `ifdef STREAM73_IN_WIDTH  | stream_in_desc_poll_next_desc[73]  `endif
                                        `ifdef STREAM73_OUT_WIDTH | stream_out_desc_poll_next_desc[73] `endif
                                        `ifdef STREAM74_IN_WIDTH  | stream_in_desc_poll_next_desc[74]  `endif
                                        `ifdef STREAM74_OUT_WIDTH | stream_out_desc_poll_next_desc[74] `endif
                                        `ifdef STREAM75_IN_WIDTH  | stream_in_desc_poll_next_desc[75]  `endif
                                        `ifdef STREAM75_OUT_WIDTH | stream_out_desc_poll_next_desc[75] `endif
                                        `ifdef STREAM76_IN_WIDTH  | stream_in_desc_poll_next_desc[76]  `endif
                                        `ifdef STREAM76_OUT_WIDTH | stream_out_desc_poll_next_desc[76] `endif
                                        `ifdef STREAM77_IN_WIDTH  | stream_in_desc_poll_next_desc[77]  `endif
                                        `ifdef STREAM77_OUT_WIDTH | stream_out_desc_poll_next_desc[77] `endif
                                        `ifdef STREAM78_IN_WIDTH  | stream_in_desc_poll_next_desc[78]  `endif
                                        `ifdef STREAM78_OUT_WIDTH | stream_out_desc_poll_next_desc[78] `endif
                                        `ifdef STREAM79_IN_WIDTH  | stream_in_desc_poll_next_desc[79]  `endif
                                        `ifdef STREAM79_OUT_WIDTH | stream_out_desc_poll_next_desc[79] `endif
                                        `ifdef STREAM80_IN_WIDTH  | stream_in_desc_poll_next_desc[80]  `endif
                                        `ifdef STREAM80_OUT_WIDTH | stream_out_desc_poll_next_desc[80] `endif
                                        `ifdef STREAM81_IN_WIDTH  | stream_in_desc_poll_next_desc[81]  `endif
                                        `ifdef STREAM81_OUT_WIDTH | stream_out_desc_poll_next_desc[81] `endif
                                        `ifdef STREAM82_IN_WIDTH  | stream_in_desc_poll_next_desc[82]  `endif
                                        `ifdef STREAM82_OUT_WIDTH | stream_out_desc_poll_next_desc[82] `endif
                                        `ifdef STREAM83_IN_WIDTH  | stream_in_desc_poll_next_desc[83]  `endif
                                        `ifdef STREAM83_OUT_WIDTH | stream_out_desc_poll_next_desc[83] `endif
                                        `ifdef STREAM84_IN_WIDTH  | stream_in_desc_poll_next_desc[84]  `endif
                                        `ifdef STREAM84_OUT_WIDTH | stream_out_desc_poll_next_desc[84] `endif
                                        `ifdef STREAM85_IN_WIDTH  | stream_in_desc_poll_next_desc[85]  `endif
                                        `ifdef STREAM85_OUT_WIDTH | stream_out_desc_poll_next_desc[85] `endif
                                        `ifdef STREAM86_IN_WIDTH  | stream_in_desc_poll_next_desc[86]  `endif
                                        `ifdef STREAM86_OUT_WIDTH | stream_out_desc_poll_next_desc[86] `endif
                                        `ifdef STREAM87_IN_WIDTH  | stream_in_desc_poll_next_desc[87]  `endif
                                        `ifdef STREAM87_OUT_WIDTH | stream_out_desc_poll_next_desc[87] `endif
                                        `ifdef STREAM88_IN_WIDTH  | stream_in_desc_poll_next_desc[88]  `endif
                                        `ifdef STREAM88_OUT_WIDTH | stream_out_desc_poll_next_desc[88] `endif
                                        `ifdef STREAM89_IN_WIDTH  | stream_in_desc_poll_next_desc[89]  `endif
                                        `ifdef STREAM89_OUT_WIDTH | stream_out_desc_poll_next_desc[89] `endif
                                        `ifdef STREAM90_IN_WIDTH  | stream_in_desc_poll_next_desc[90]  `endif
                                        `ifdef STREAM90_OUT_WIDTH | stream_out_desc_poll_next_desc[90] `endif
                                        `ifdef STREAM91_IN_WIDTH  | stream_in_desc_poll_next_desc[91]  `endif
                                        `ifdef STREAM91_OUT_WIDTH | stream_out_desc_poll_next_desc[91] `endif
                                        `ifdef STREAM92_IN_WIDTH  | stream_in_desc_poll_next_desc[92]  `endif
                                        `ifdef STREAM92_OUT_WIDTH | stream_out_desc_poll_next_desc[92] `endif
                                        `ifdef STREAM93_IN_WIDTH  | stream_in_desc_poll_next_desc[93]  `endif
                                        `ifdef STREAM93_OUT_WIDTH | stream_out_desc_poll_next_desc[93] `endif
                                        `ifdef STREAM94_IN_WIDTH  | stream_in_desc_poll_next_desc[94]  `endif
                                        `ifdef STREAM94_OUT_WIDTH | stream_out_desc_poll_next_desc[94] `endif
                                        `ifdef STREAM95_IN_WIDTH  | stream_in_desc_poll_next_desc[95]  `endif
                                        `ifdef STREAM95_OUT_WIDTH | stream_out_desc_poll_next_desc[95] `endif
                                        `ifdef STREAM96_IN_WIDTH  | stream_in_desc_poll_next_desc[96]  `endif
                                        `ifdef STREAM96_OUT_WIDTH | stream_out_desc_poll_next_desc[96] `endif
                                        `ifdef STREAM97_IN_WIDTH  | stream_in_desc_poll_next_desc[97]  `endif
                                        `ifdef STREAM97_OUT_WIDTH | stream_out_desc_poll_next_desc[97] `endif
                                        `ifdef STREAM98_IN_WIDTH  | stream_in_desc_poll_next_desc[98]  `endif
                                        `ifdef STREAM98_OUT_WIDTH | stream_out_desc_poll_next_desc[98] `endif
                                        `ifdef STREAM99_IN_WIDTH  | stream_in_desc_poll_next_desc[99]  `endif
                                        `ifdef STREAM99_OUT_WIDTH | stream_out_desc_poll_next_desc[99] `endif
                                        `ifdef STREAM100_IN_WIDTH  | stream_in_desc_poll_next_desc[100]  `endif
                                        `ifdef STREAM100_OUT_WIDTH | stream_out_desc_poll_next_desc[100] `endif
                                        `ifdef STREAM101_IN_WIDTH  | stream_in_desc_poll_next_desc[101]  `endif
                                        `ifdef STREAM101_OUT_WIDTH | stream_out_desc_poll_next_desc[101] `endif
                                        `ifdef STREAM102_IN_WIDTH  | stream_in_desc_poll_next_desc[102]  `endif
                                        `ifdef STREAM102_OUT_WIDTH | stream_out_desc_poll_next_desc[102] `endif
                                        `ifdef STREAM103_IN_WIDTH  | stream_in_desc_poll_next_desc[103]  `endif
                                        `ifdef STREAM103_OUT_WIDTH | stream_out_desc_poll_next_desc[103] `endif
                                        `ifdef STREAM104_IN_WIDTH  | stream_in_desc_poll_next_desc[104]  `endif
                                        `ifdef STREAM104_OUT_WIDTH | stream_out_desc_poll_next_desc[104] `endif
                                        `ifdef STREAM105_IN_WIDTH  | stream_in_desc_poll_next_desc[105]  `endif
                                        `ifdef STREAM105_OUT_WIDTH | stream_out_desc_poll_next_desc[105] `endif
                                        `ifdef STREAM106_IN_WIDTH  | stream_in_desc_poll_next_desc[106]  `endif
                                        `ifdef STREAM106_OUT_WIDTH | stream_out_desc_poll_next_desc[106] `endif
                                        `ifdef STREAM107_IN_WIDTH  | stream_in_desc_poll_next_desc[107]  `endif
                                        `ifdef STREAM107_OUT_WIDTH | stream_out_desc_poll_next_desc[107] `endif
                                        `ifdef STREAM108_IN_WIDTH  | stream_in_desc_poll_next_desc[108]  `endif
                                        `ifdef STREAM108_OUT_WIDTH | stream_out_desc_poll_next_desc[108] `endif
                                        `ifdef STREAM109_IN_WIDTH  | stream_in_desc_poll_next_desc[109]  `endif
                                        `ifdef STREAM109_OUT_WIDTH | stream_out_desc_poll_next_desc[109] `endif
                                        `ifdef STREAM110_IN_WIDTH  | stream_in_desc_poll_next_desc[110]  `endif
                                        `ifdef STREAM110_OUT_WIDTH | stream_out_desc_poll_next_desc[110] `endif
                                        `ifdef STREAM111_IN_WIDTH  | stream_in_desc_poll_next_desc[111]  `endif
                                        `ifdef STREAM111_OUT_WIDTH | stream_out_desc_poll_next_desc[111] `endif
                                        `ifdef STREAM112_IN_WIDTH  | stream_in_desc_poll_next_desc[112]  `endif
                                        `ifdef STREAM112_OUT_WIDTH | stream_out_desc_poll_next_desc[112] `endif
                                        `ifdef STREAM113_IN_WIDTH  | stream_in_desc_poll_next_desc[113]  `endif
                                        `ifdef STREAM113_OUT_WIDTH | stream_out_desc_poll_next_desc[113] `endif
                                        `ifdef STREAM114_IN_WIDTH  | stream_in_desc_poll_next_desc[114]  `endif
                                        `ifdef STREAM114_OUT_WIDTH | stream_out_desc_poll_next_desc[114] `endif
                                        `ifdef STREAM115_IN_WIDTH  | stream_in_desc_poll_next_desc[115]  `endif
                                        `ifdef STREAM115_OUT_WIDTH | stream_out_desc_poll_next_desc[115] `endif
                                        `ifdef STREAM116_IN_WIDTH  | stream_in_desc_poll_next_desc[116]  `endif
                                        `ifdef STREAM116_OUT_WIDTH | stream_out_desc_poll_next_desc[116] `endif
                                        `ifdef STREAM117_IN_WIDTH  | stream_in_desc_poll_next_desc[117]  `endif
                                        `ifdef STREAM117_OUT_WIDTH | stream_out_desc_poll_next_desc[117] `endif
                                        `ifdef STREAM118_IN_WIDTH  | stream_in_desc_poll_next_desc[118]  `endif
                                        `ifdef STREAM118_OUT_WIDTH | stream_out_desc_poll_next_desc[118] `endif
                                        `ifdef STREAM119_IN_WIDTH  | stream_in_desc_poll_next_desc[119]  `endif
                                        `ifdef STREAM119_OUT_WIDTH | stream_out_desc_poll_next_desc[119] `endif
                                        `ifdef STREAM120_IN_WIDTH  | stream_in_desc_poll_next_desc[120]  `endif
                                        `ifdef STREAM120_OUT_WIDTH | stream_out_desc_poll_next_desc[120] `endif
                                        `ifdef STREAM121_IN_WIDTH  | stream_in_desc_poll_next_desc[121]  `endif
                                        `ifdef STREAM121_OUT_WIDTH | stream_out_desc_poll_next_desc[121] `endif
                                        `ifdef STREAM122_IN_WIDTH  | stream_in_desc_poll_next_desc[122]  `endif
                                        `ifdef STREAM122_OUT_WIDTH | stream_out_desc_poll_next_desc[122] `endif
                                        `ifdef STREAM123_IN_WIDTH  | stream_in_desc_poll_next_desc[123]  `endif
                                        `ifdef STREAM123_OUT_WIDTH | stream_out_desc_poll_next_desc[123] `endif
                                        `ifdef STREAM124_IN_WIDTH  | stream_in_desc_poll_next_desc[124]  `endif
                                        `ifdef STREAM124_OUT_WIDTH | stream_out_desc_poll_next_desc[124] `endif
                                        `ifdef STREAM125_IN_WIDTH  | stream_in_desc_poll_next_desc[125]  `endif
                                        `ifdef STREAM125_OUT_WIDTH | stream_out_desc_poll_next_desc[125] `endif
                                        `ifdef STREAM126_IN_WIDTH  | stream_in_desc_poll_next_desc[126]  `endif
                                        `ifdef STREAM126_OUT_WIDTH | stream_out_desc_poll_next_desc[126] `endif
                                        );
    assign s_out_data[C_DATA_WIDTH-1:0] = ({C_DATA_WIDTH{1'b0}}
                                        `ifdef PICOBUS_WIDTH | s_out_data_userpb `endif
                                        `ifdef STREAM1_OUT_WIDTH | stream_out_data_card[1][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM2_OUT_WIDTH | stream_out_data_card[2][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM3_OUT_WIDTH | stream_out_data_card[3][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM4_OUT_WIDTH | stream_out_data_card[4][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM5_OUT_WIDTH | stream_out_data_card[5][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM6_OUT_WIDTH | stream_out_data_card[6][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM7_OUT_WIDTH | stream_out_data_card[7][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM8_OUT_WIDTH | stream_out_data_card[8][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM9_OUT_WIDTH | stream_out_data_card[9][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM10_OUT_WIDTH | stream_out_data_card[10][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM11_OUT_WIDTH | stream_out_data_card[11][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM12_OUT_WIDTH | stream_out_data_card[12][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM13_OUT_WIDTH | stream_out_data_card[13][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM14_OUT_WIDTH | stream_out_data_card[14][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM15_OUT_WIDTH | stream_out_data_card[15][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM16_OUT_WIDTH | stream_out_data_card[16][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM17_OUT_WIDTH | stream_out_data_card[17][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM18_OUT_WIDTH | stream_out_data_card[18][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM19_OUT_WIDTH | stream_out_data_card[19][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM20_OUT_WIDTH | stream_out_data_card[20][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM21_OUT_WIDTH | stream_out_data_card[21][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM22_OUT_WIDTH | stream_out_data_card[22][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM23_OUT_WIDTH | stream_out_data_card[23][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM24_OUT_WIDTH | stream_out_data_card[24][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM25_OUT_WIDTH | stream_out_data_card[25][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM26_OUT_WIDTH | stream_out_data_card[26][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM27_OUT_WIDTH | stream_out_data_card[27][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM28_OUT_WIDTH | stream_out_data_card[28][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM29_OUT_WIDTH | stream_out_data_card[29][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM30_OUT_WIDTH | stream_out_data_card[30][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM31_OUT_WIDTH | stream_out_data_card[31][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM32_OUT_WIDTH | stream_out_data_card[32][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM33_OUT_WIDTH | stream_out_data_card[33][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM34_OUT_WIDTH | stream_out_data_card[34][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM35_OUT_WIDTH | stream_out_data_card[35][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM36_OUT_WIDTH | stream_out_data_card[36][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM37_OUT_WIDTH | stream_out_data_card[37][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM38_OUT_WIDTH | stream_out_data_card[38][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM39_OUT_WIDTH | stream_out_data_card[39][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM40_OUT_WIDTH | stream_out_data_card[40][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM41_OUT_WIDTH | stream_out_data_card[41][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM42_OUT_WIDTH | stream_out_data_card[42][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM43_OUT_WIDTH | stream_out_data_card[43][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM44_OUT_WIDTH | stream_out_data_card[44][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM45_OUT_WIDTH | stream_out_data_card[45][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM46_OUT_WIDTH | stream_out_data_card[46][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM47_OUT_WIDTH | stream_out_data_card[47][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM48_OUT_WIDTH | stream_out_data_card[48][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM49_OUT_WIDTH | stream_out_data_card[49][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM50_OUT_WIDTH | stream_out_data_card[50][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM51_OUT_WIDTH | stream_out_data_card[51][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM52_OUT_WIDTH | stream_out_data_card[52][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM53_OUT_WIDTH | stream_out_data_card[53][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM54_OUT_WIDTH | stream_out_data_card[54][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM55_OUT_WIDTH | stream_out_data_card[55][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM56_OUT_WIDTH | stream_out_data_card[56][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM57_OUT_WIDTH | stream_out_data_card[57][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM58_OUT_WIDTH | stream_out_data_card[58][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM59_OUT_WIDTH | stream_out_data_card[59][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM60_OUT_WIDTH | stream_out_data_card[60][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM61_OUT_WIDTH | stream_out_data_card[61][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM62_OUT_WIDTH | stream_out_data_card[62][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM63_OUT_WIDTH | stream_out_data_card[63][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM64_OUT_WIDTH | stream_out_data_card[64][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM65_OUT_WIDTH | stream_out_data_card[65][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM66_OUT_WIDTH | stream_out_data_card[66][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM67_OUT_WIDTH | stream_out_data_card[67][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM68_OUT_WIDTH | stream_out_data_card[68][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM69_OUT_WIDTH | stream_out_data_card[69][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM70_OUT_WIDTH | stream_out_data_card[70][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM71_OUT_WIDTH | stream_out_data_card[71][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM72_OUT_WIDTH | stream_out_data_card[72][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM73_OUT_WIDTH | stream_out_data_card[73][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM74_OUT_WIDTH | stream_out_data_card[74][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM75_OUT_WIDTH | stream_out_data_card[75][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM76_OUT_WIDTH | stream_out_data_card[76][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM77_OUT_WIDTH | stream_out_data_card[77][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM78_OUT_WIDTH | stream_out_data_card[78][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM79_OUT_WIDTH | stream_out_data_card[79][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM80_OUT_WIDTH | stream_out_data_card[80][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM81_OUT_WIDTH | stream_out_data_card[81][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM82_OUT_WIDTH | stream_out_data_card[82][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM83_OUT_WIDTH | stream_out_data_card[83][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM84_OUT_WIDTH | stream_out_data_card[84][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM85_OUT_WIDTH | stream_out_data_card[85][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM86_OUT_WIDTH | stream_out_data_card[86][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM87_OUT_WIDTH | stream_out_data_card[87][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM88_OUT_WIDTH | stream_out_data_card[88][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM89_OUT_WIDTH | stream_out_data_card[89][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM90_OUT_WIDTH | stream_out_data_card[90][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM91_OUT_WIDTH | stream_out_data_card[91][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM92_OUT_WIDTH | stream_out_data_card[92][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM93_OUT_WIDTH | stream_out_data_card[93][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM94_OUT_WIDTH | stream_out_data_card[94][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM95_OUT_WIDTH | stream_out_data_card[95][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM96_OUT_WIDTH | stream_out_data_card[96][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM97_OUT_WIDTH | stream_out_data_card[97][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM98_OUT_WIDTH | stream_out_data_card[98][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM99_OUT_WIDTH | stream_out_data_card[99][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM100_OUT_WIDTH | stream_out_data_card[100][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM101_OUT_WIDTH | stream_out_data_card[101][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM102_OUT_WIDTH | stream_out_data_card[102][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM103_OUT_WIDTH | stream_out_data_card[103][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM104_OUT_WIDTH | stream_out_data_card[104][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM105_OUT_WIDTH | stream_out_data_card[105][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM106_OUT_WIDTH | stream_out_data_card[106][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM107_OUT_WIDTH | stream_out_data_card[107][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM108_OUT_WIDTH | stream_out_data_card[108][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM109_OUT_WIDTH | stream_out_data_card[109][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM110_OUT_WIDTH | stream_out_data_card[110][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM111_OUT_WIDTH | stream_out_data_card[111][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM112_OUT_WIDTH | stream_out_data_card[112][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM113_OUT_WIDTH | stream_out_data_card[113][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM114_OUT_WIDTH | stream_out_data_card[114][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM115_OUT_WIDTH | stream_out_data_card[115][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM116_OUT_WIDTH | stream_out_data_card[116][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM117_OUT_WIDTH | stream_out_data_card[117][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM118_OUT_WIDTH | stream_out_data_card[118][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM119_OUT_WIDTH | stream_out_data_card[119][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM120_OUT_WIDTH | stream_out_data_card[120][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM121_OUT_WIDTH | stream_out_data_card[121][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM122_OUT_WIDTH | stream_out_data_card[122][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM123_OUT_WIDTH | stream_out_data_card[123][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM124_OUT_WIDTH | stream_out_data_card[124][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM125_OUT_WIDTH | stream_out_data_card[125][C_DATA_WIDTH-1:0] `endif
                                        `ifdef STREAM126_OUT_WIDTH | stream_out_data_card[126][C_DATA_WIDTH-1:0] `endif
                                        );
    assign s_out_ow_dvld[OW_DVLD_W-1:0] = ({OW_DVLD_W{1'b0}}
                                        `ifdef PICOBUS_WIDTH | s_out_ow_dvld_userpb `endif
                                        `ifdef STREAM1_OUT_WIDTH | stream_out_ow_dvld_card[1][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM2_OUT_WIDTH | stream_out_ow_dvld_card[2][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM3_OUT_WIDTH | stream_out_ow_dvld_card[3][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM4_OUT_WIDTH | stream_out_ow_dvld_card[4][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM5_OUT_WIDTH | stream_out_ow_dvld_card[5][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM6_OUT_WIDTH | stream_out_ow_dvld_card[6][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM7_OUT_WIDTH | stream_out_ow_dvld_card[7][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM8_OUT_WIDTH | stream_out_ow_dvld_card[8][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM9_OUT_WIDTH | stream_out_ow_dvld_card[9][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM10_OUT_WIDTH | stream_out_ow_dvld_card[10][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM11_OUT_WIDTH | stream_out_ow_dvld_card[11][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM12_OUT_WIDTH | stream_out_ow_dvld_card[12][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM13_OUT_WIDTH | stream_out_ow_dvld_card[13][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM14_OUT_WIDTH | stream_out_ow_dvld_card[14][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM15_OUT_WIDTH | stream_out_ow_dvld_card[15][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM16_OUT_WIDTH | stream_out_ow_dvld_card[16][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM17_OUT_WIDTH | stream_out_ow_dvld_card[17][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM18_OUT_WIDTH | stream_out_ow_dvld_card[18][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM19_OUT_WIDTH | stream_out_ow_dvld_card[19][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM20_OUT_WIDTH | stream_out_ow_dvld_card[20][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM21_OUT_WIDTH | stream_out_ow_dvld_card[21][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM22_OUT_WIDTH | stream_out_ow_dvld_card[22][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM23_OUT_WIDTH | stream_out_ow_dvld_card[23][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM24_OUT_WIDTH | stream_out_ow_dvld_card[24][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM25_OUT_WIDTH | stream_out_ow_dvld_card[25][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM26_OUT_WIDTH | stream_out_ow_dvld_card[26][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM27_OUT_WIDTH | stream_out_ow_dvld_card[27][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM28_OUT_WIDTH | stream_out_ow_dvld_card[28][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM29_OUT_WIDTH | stream_out_ow_dvld_card[29][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM30_OUT_WIDTH | stream_out_ow_dvld_card[30][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM31_OUT_WIDTH | stream_out_ow_dvld_card[31][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM32_OUT_WIDTH | stream_out_ow_dvld_card[32][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM33_OUT_WIDTH | stream_out_ow_dvld_card[33][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM34_OUT_WIDTH | stream_out_ow_dvld_card[34][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM35_OUT_WIDTH | stream_out_ow_dvld_card[35][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM36_OUT_WIDTH | stream_out_ow_dvld_card[36][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM37_OUT_WIDTH | stream_out_ow_dvld_card[37][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM38_OUT_WIDTH | stream_out_ow_dvld_card[38][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM39_OUT_WIDTH | stream_out_ow_dvld_card[39][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM40_OUT_WIDTH | stream_out_ow_dvld_card[40][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM41_OUT_WIDTH | stream_out_ow_dvld_card[41][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM42_OUT_WIDTH | stream_out_ow_dvld_card[42][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM43_OUT_WIDTH | stream_out_ow_dvld_card[43][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM44_OUT_WIDTH | stream_out_ow_dvld_card[44][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM45_OUT_WIDTH | stream_out_ow_dvld_card[45][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM46_OUT_WIDTH | stream_out_ow_dvld_card[46][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM47_OUT_WIDTH | stream_out_ow_dvld_card[47][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM48_OUT_WIDTH | stream_out_ow_dvld_card[48][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM49_OUT_WIDTH | stream_out_ow_dvld_card[49][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM50_OUT_WIDTH | stream_out_ow_dvld_card[50][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM51_OUT_WIDTH | stream_out_ow_dvld_card[51][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM52_OUT_WIDTH | stream_out_ow_dvld_card[52][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM53_OUT_WIDTH | stream_out_ow_dvld_card[53][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM54_OUT_WIDTH | stream_out_ow_dvld_card[54][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM55_OUT_WIDTH | stream_out_ow_dvld_card[55][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM56_OUT_WIDTH | stream_out_ow_dvld_card[56][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM57_OUT_WIDTH | stream_out_ow_dvld_card[57][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM58_OUT_WIDTH | stream_out_ow_dvld_card[58][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM59_OUT_WIDTH | stream_out_ow_dvld_card[59][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM60_OUT_WIDTH | stream_out_ow_dvld_card[60][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM61_OUT_WIDTH | stream_out_ow_dvld_card[61][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM62_OUT_WIDTH | stream_out_ow_dvld_card[62][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM63_OUT_WIDTH | stream_out_ow_dvld_card[63][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM64_OUT_WIDTH | stream_out_ow_dvld_card[64][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM65_OUT_WIDTH | stream_out_ow_dvld_card[65][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM66_OUT_WIDTH | stream_out_ow_dvld_card[66][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM67_OUT_WIDTH | stream_out_ow_dvld_card[67][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM68_OUT_WIDTH | stream_out_ow_dvld_card[68][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM69_OUT_WIDTH | stream_out_ow_dvld_card[69][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM70_OUT_WIDTH | stream_out_ow_dvld_card[70][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM71_OUT_WIDTH | stream_out_ow_dvld_card[71][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM72_OUT_WIDTH | stream_out_ow_dvld_card[72][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM73_OUT_WIDTH | stream_out_ow_dvld_card[73][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM74_OUT_WIDTH | stream_out_ow_dvld_card[74][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM75_OUT_WIDTH | stream_out_ow_dvld_card[75][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM76_OUT_WIDTH | stream_out_ow_dvld_card[76][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM77_OUT_WIDTH | stream_out_ow_dvld_card[77][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM78_OUT_WIDTH | stream_out_ow_dvld_card[78][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM79_OUT_WIDTH | stream_out_ow_dvld_card[79][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM80_OUT_WIDTH | stream_out_ow_dvld_card[80][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM81_OUT_WIDTH | stream_out_ow_dvld_card[81][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM82_OUT_WIDTH | stream_out_ow_dvld_card[82][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM83_OUT_WIDTH | stream_out_ow_dvld_card[83][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM84_OUT_WIDTH | stream_out_ow_dvld_card[84][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM85_OUT_WIDTH | stream_out_ow_dvld_card[85][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM86_OUT_WIDTH | stream_out_ow_dvld_card[86][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM87_OUT_WIDTH | stream_out_ow_dvld_card[87][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM88_OUT_WIDTH | stream_out_ow_dvld_card[88][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM89_OUT_WIDTH | stream_out_ow_dvld_card[89][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM90_OUT_WIDTH | stream_out_ow_dvld_card[90][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM91_OUT_WIDTH | stream_out_ow_dvld_card[91][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM92_OUT_WIDTH | stream_out_ow_dvld_card[92][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM93_OUT_WIDTH | stream_out_ow_dvld_card[93][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM94_OUT_WIDTH | stream_out_ow_dvld_card[94][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM95_OUT_WIDTH | stream_out_ow_dvld_card[95][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM96_OUT_WIDTH | stream_out_ow_dvld_card[96][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM97_OUT_WIDTH | stream_out_ow_dvld_card[97][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM98_OUT_WIDTH | stream_out_ow_dvld_card[98][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM99_OUT_WIDTH | stream_out_ow_dvld_card[99][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM100_OUT_WIDTH | stream_out_ow_dvld_card[100][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM101_OUT_WIDTH | stream_out_ow_dvld_card[101][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM102_OUT_WIDTH | stream_out_ow_dvld_card[102][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM103_OUT_WIDTH | stream_out_ow_dvld_card[103][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM104_OUT_WIDTH | stream_out_ow_dvld_card[104][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM105_OUT_WIDTH | stream_out_ow_dvld_card[105][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM106_OUT_WIDTH | stream_out_ow_dvld_card[106][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM107_OUT_WIDTH | stream_out_ow_dvld_card[107][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM108_OUT_WIDTH | stream_out_ow_dvld_card[108][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM109_OUT_WIDTH | stream_out_ow_dvld_card[109][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM110_OUT_WIDTH | stream_out_ow_dvld_card[110][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM111_OUT_WIDTH | stream_out_ow_dvld_card[111][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM112_OUT_WIDTH | stream_out_ow_dvld_card[112][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM113_OUT_WIDTH | stream_out_ow_dvld_card[113][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM114_OUT_WIDTH | stream_out_ow_dvld_card[114][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM115_OUT_WIDTH | stream_out_ow_dvld_card[115][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM116_OUT_WIDTH | stream_out_ow_dvld_card[116][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM117_OUT_WIDTH | stream_out_ow_dvld_card[117][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM118_OUT_WIDTH | stream_out_ow_dvld_card[118][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM119_OUT_WIDTH | stream_out_ow_dvld_card[119][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM120_OUT_WIDTH | stream_out_ow_dvld_card[120][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM121_OUT_WIDTH | stream_out_ow_dvld_card[121][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM122_OUT_WIDTH | stream_out_ow_dvld_card[122][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM123_OUT_WIDTH | stream_out_ow_dvld_card[123][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM124_OUT_WIDTH | stream_out_ow_dvld_card[124][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM125_OUT_WIDTH | stream_out_ow_dvld_card[125][OW_DVLD_W-1:0] `endif
                                        `ifdef STREAM126_OUT_WIDTH | stream_out_ow_dvld_card[126][OW_DVLD_W-1:0] `endif
                                        );


endmodule

